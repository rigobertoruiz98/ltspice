* C:\Users\ruizc\Downloads\knowles\knowles.asc
m:x1:1 vdd x1:na x1:n001 vdd x1:pfet l=0.6u w=6u
m:x1:2 x1:n001 b1 p1 vdd x1:pfet l=0.6u w=6u
m:x1:3 vdd a1 x1:n002 vdd x1:pfet l=0.6u w=6u
m:x1:4 x1:n002 x1:nb p1 vdd x1:pfet l=0.6u w=6u
m:x1:5 p1 b1 x1:n004 0 x1:nfet l=0.6u w=3u
m:x1:6 x1:n004 a1 0 0 x1:nfet l=0.6u w=3u
m:x1:7 p1 x1:nb x1:n005 0 x1:nfet l=0.6u w=3u
m:x1:8 x1:n005 x1:na 0 0 x1:nfet l=0.6u w=3u
m:x1:9 vdd b1 x1:nb vdd x1:pfet l=0.6u w=3u
m:x1:10 x1:nb b1 0 0 x1:nfet l=0.6u w=1.5u
m:x1:11 vdd a1 x1:na vdd x1:pfet l=0.6u w=3u
m:x1:12 x1:na a1 0 0 x1:nfet l=0.6u w=1.5u
m:x1:13 x1:nand b1 x1:n003 0 x1:nfet l=0.6u w=3u
m:x1:14 x1:n003 a1 0 0 x1:nfet l=0.6u w=3u
m:x1:15 vdd a1 x1:nand vdd x1:pfet l=0.6u w=3u
m:x1:16 vdd b1 x1:nand vdd x1:pfet l=0.6u w=3u
m:x1:17 vdd x1:nand n014 vdd x1:pfet l=0.6u w=3u
m:x1:18 n014 x1:nand 0 0 x1:nfet l=0.6u w=1.5u
m:x2:1 vdd x2:na x2:n001 vdd x2:pfet l=0.6u w=6u
m:x2:2 x2:n001 b2 p2 vdd x2:pfet l=0.6u w=6u
m:x2:3 vdd a2 x2:n002 vdd x2:pfet l=0.6u w=6u
m:x2:4 x2:n002 x2:nb p2 vdd x2:pfet l=0.6u w=6u
m:x2:5 p2 b2 x2:n004 0 x2:nfet l=0.6u w=3u
m:x2:6 x2:n004 a2 0 0 x2:nfet l=0.6u w=3u
m:x2:7 p2 x2:nb x2:n005 0 x2:nfet l=0.6u w=3u
m:x2:8 x2:n005 x2:na 0 0 x2:nfet l=0.6u w=3u
m:x2:9 vdd b2 x2:nb vdd x2:pfet l=0.6u w=3u
m:x2:10 x2:nb b2 0 0 x2:nfet l=0.6u w=1.5u
m:x2:11 vdd a2 x2:na vdd x2:pfet l=0.6u w=3u
m:x2:12 x2:na a2 0 0 x2:nfet l=0.6u w=1.5u
m:x2:13 x2:nand b2 x2:n003 0 x2:nfet l=0.6u w=3u
m:x2:14 x2:n003 a2 0 0 x2:nfet l=0.6u w=3u
m:x2:15 vdd a2 x2:nand vdd x2:pfet l=0.6u w=3u
m:x2:16 vdd b2 x2:nand vdd x2:pfet l=0.6u w=3u
m:x2:17 vdd x2:nand n013 vdd x2:pfet l=0.6u w=3u
m:x2:18 n013 x2:nand 0 0 x2:nfet l=0.6u w=1.5u
m:x3:1 vdd x3:na x3:n001 vdd x3:pfet l=0.6u w=6u
m:x3:2 x3:n001 b3 p3 vdd x3:pfet l=0.6u w=6u
m:x3:3 vdd a3 x3:n002 vdd x3:pfet l=0.6u w=6u
m:x3:4 x3:n002 x3:nb p3 vdd x3:pfet l=0.6u w=6u
m:x3:5 p3 b3 x3:n004 0 x3:nfet l=0.6u w=3u
m:x3:6 x3:n004 a3 0 0 x3:nfet l=0.6u w=3u
m:x3:7 p3 x3:nb x3:n005 0 x3:nfet l=0.6u w=3u
m:x3:8 x3:n005 x3:na 0 0 x3:nfet l=0.6u w=3u
m:x3:9 vdd b3 x3:nb vdd x3:pfet l=0.6u w=3u
m:x3:10 x3:nb b3 0 0 x3:nfet l=0.6u w=1.5u
m:x3:11 vdd a3 x3:na vdd x3:pfet l=0.6u w=3u
m:x3:12 x3:na a3 0 0 x3:nfet l=0.6u w=1.5u
m:x3:13 x3:nand b3 x3:n003 0 x3:nfet l=0.6u w=3u
m:x3:14 x3:n003 a3 0 0 x3:nfet l=0.6u w=3u
m:x3:15 vdd a3 x3:nand vdd x3:pfet l=0.6u w=3u
m:x3:16 vdd b3 x3:nand vdd x3:pfet l=0.6u w=3u
m:x3:17 vdd x3:nand n012 vdd x3:pfet l=0.6u w=3u
m:x3:18 n012 x3:nand 0 0 x3:nfet l=0.6u w=1.5u
m:x4:1 vdd x4:na x4:n001 vdd x4:pfet l=0.6u w=6u
m:x4:2 x4:n001 b4 p4 vdd x4:pfet l=0.6u w=6u
m:x4:3 vdd a4 x4:n002 vdd x4:pfet l=0.6u w=6u
m:x4:4 x4:n002 x4:nb p4 vdd x4:pfet l=0.6u w=6u
m:x4:5 p4 b4 x4:n004 0 x4:nfet l=0.6u w=3u
m:x4:6 x4:n004 a4 0 0 x4:nfet l=0.6u w=3u
m:x4:7 p4 x4:nb x4:n005 0 x4:nfet l=0.6u w=3u
m:x4:8 x4:n005 x4:na 0 0 x4:nfet l=0.6u w=3u
m:x4:9 vdd b4 x4:nb vdd x4:pfet l=0.6u w=3u
m:x4:10 x4:nb b4 0 0 x4:nfet l=0.6u w=1.5u
m:x4:11 vdd a4 x4:na vdd x4:pfet l=0.6u w=3u
m:x4:12 x4:na a4 0 0 x4:nfet l=0.6u w=1.5u
m:x4:13 x4:nand b4 x4:n003 0 x4:nfet l=0.6u w=3u
m:x4:14 x4:n003 a4 0 0 x4:nfet l=0.6u w=3u
m:x4:15 vdd a4 x4:nand vdd x4:pfet l=0.6u w=3u
m:x4:16 vdd b4 x4:nand vdd x4:pfet l=0.6u w=3u
m:x4:17 vdd x4:nand n011 vdd x4:pfet l=0.6u w=3u
m:x4:18 n011 x4:nand 0 0 x4:nfet l=0.6u w=1.5u
m:x5:1 vdd x5:na x5:n001 vdd x5:pfet l=0.6u w=6u
m:x5:2 x5:n001 b5 p5 vdd x5:pfet l=0.6u w=6u
m:x5:3 vdd a5 x5:n002 vdd x5:pfet l=0.6u w=6u
m:x5:4 x5:n002 x5:nb p5 vdd x5:pfet l=0.6u w=6u
m:x5:5 p5 b5 x5:n004 0 x5:nfet l=0.6u w=3u
m:x5:6 x5:n004 a5 0 0 x5:nfet l=0.6u w=3u
m:x5:7 p5 x5:nb x5:n005 0 x5:nfet l=0.6u w=3u
m:x5:8 x5:n005 x5:na 0 0 x5:nfet l=0.6u w=3u
m:x5:9 vdd b5 x5:nb vdd x5:pfet l=0.6u w=3u
m:x5:10 x5:nb b5 0 0 x5:nfet l=0.6u w=1.5u
m:x5:11 vdd a5 x5:na vdd x5:pfet l=0.6u w=3u
m:x5:12 x5:na a5 0 0 x5:nfet l=0.6u w=1.5u
m:x5:13 x5:nand b5 x5:n003 0 x5:nfet l=0.6u w=3u
m:x5:14 x5:n003 a5 0 0 x5:nfet l=0.6u w=3u
m:x5:15 vdd a5 x5:nand vdd x5:pfet l=0.6u w=3u
m:x5:16 vdd b5 x5:nand vdd x5:pfet l=0.6u w=3u
m:x5:17 vdd x5:nand n010 vdd x5:pfet l=0.6u w=3u
m:x5:18 n010 x5:nand 0 0 x5:nfet l=0.6u w=1.5u
m:x6:1 vdd x6:na x6:n001 vdd x6:pfet l=0.6u w=6u
m:x6:2 x6:n001 b6 p6 vdd x6:pfet l=0.6u w=6u
m:x6:3 vdd a6 x6:n002 vdd x6:pfet l=0.6u w=6u
m:x6:4 x6:n002 x6:nb p6 vdd x6:pfet l=0.6u w=6u
m:x6:5 p6 b6 x6:n004 0 x6:nfet l=0.6u w=3u
m:x6:6 x6:n004 a6 0 0 x6:nfet l=0.6u w=3u
m:x6:7 p6 x6:nb x6:n005 0 x6:nfet l=0.6u w=3u
m:x6:8 x6:n005 x6:na 0 0 x6:nfet l=0.6u w=3u
m:x6:9 vdd b6 x6:nb vdd x6:pfet l=0.6u w=3u
m:x6:10 x6:nb b6 0 0 x6:nfet l=0.6u w=1.5u
m:x6:11 vdd a6 x6:na vdd x6:pfet l=0.6u w=3u
m:x6:12 x6:na a6 0 0 x6:nfet l=0.6u w=1.5u
m:x6:13 x6:nand b6 x6:n003 0 x6:nfet l=0.6u w=3u
m:x6:14 x6:n003 a6 0 0 x6:nfet l=0.6u w=3u
m:x6:15 vdd a6 x6:nand vdd x6:pfet l=0.6u w=3u
m:x6:16 vdd b6 x6:nand vdd x6:pfet l=0.6u w=3u
m:x6:17 vdd x6:nand n009 vdd x6:pfet l=0.6u w=3u
m:x6:18 n009 x6:nand 0 0 x6:nfet l=0.6u w=1.5u
m:x7:1 vdd x7:na x7:n001 vdd x7:pfet l=0.6u w=6u
m:x7:2 x7:n001 b7 p7 vdd x7:pfet l=0.6u w=6u
m:x7:3 vdd a7 x7:n002 vdd x7:pfet l=0.6u w=6u
m:x7:4 x7:n002 x7:nb p7 vdd x7:pfet l=0.6u w=6u
m:x7:5 p7 b7 x7:n004 0 x7:nfet l=0.6u w=3u
m:x7:6 x7:n004 a7 0 0 x7:nfet l=0.6u w=3u
m:x7:7 p7 x7:nb x7:n005 0 x7:nfet l=0.6u w=3u
m:x7:8 x7:n005 x7:na 0 0 x7:nfet l=0.6u w=3u
m:x7:9 vdd b7 x7:nb vdd x7:pfet l=0.6u w=3u
m:x7:10 x7:nb b7 0 0 x7:nfet l=0.6u w=1.5u
m:x7:11 vdd a7 x7:na vdd x7:pfet l=0.6u w=3u
m:x7:12 x7:na a7 0 0 x7:nfet l=0.6u w=1.5u
m:x7:13 x7:nand b7 x7:n003 0 x7:nfet l=0.6u w=3u
m:x7:14 x7:n003 a7 0 0 x7:nfet l=0.6u w=3u
m:x7:15 vdd a7 x7:nand vdd x7:pfet l=0.6u w=3u
m:x7:16 vdd b7 x7:nand vdd x7:pfet l=0.6u w=3u
m:x7:17 vdd x7:nand n008 vdd x7:pfet l=0.6u w=3u
m:x7:18 n008 x7:nand 0 0 x7:nfet l=0.6u w=1.5u
m:x8:1 vdd x8:na x8:n001 vdd x8:pfet l=0.6u w=6u
m:x8:2 x8:n001 b8 p8 vdd x8:pfet l=0.6u w=6u
m:x8:3 vdd a8 x8:n002 vdd x8:pfet l=0.6u w=6u
m:x8:4 x8:n002 x8:nb p8 vdd x8:pfet l=0.6u w=6u
m:x8:5 p8 b8 x8:n004 0 x8:nfet l=0.6u w=3u
m:x8:6 x8:n004 a8 0 0 x8:nfet l=0.6u w=3u
m:x8:7 p8 x8:nb x8:n005 0 x8:nfet l=0.6u w=3u
m:x8:8 x8:n005 x8:na 0 0 x8:nfet l=0.6u w=3u
m:x8:9 vdd b8 x8:nb vdd x8:pfet l=0.6u w=3u
m:x8:10 x8:nb b8 0 0 x8:nfet l=0.6u w=1.5u
m:x8:11 vdd a8 x8:na vdd x8:pfet l=0.6u w=3u
m:x8:12 x8:na a8 0 0 x8:nfet l=0.6u w=1.5u
m:x8:13 x8:nand b8 x8:n003 0 x8:nfet l=0.6u w=3u
m:x8:14 x8:n003 a8 0 0 x8:nfet l=0.6u w=3u
m:x8:15 vdd a8 x8:nand vdd x8:pfet l=0.6u w=3u
m:x8:16 vdd b8 x8:nand vdd x8:pfet l=0.6u w=3u
m:x8:17 vdd x8:nand n007 vdd x8:pfet l=0.6u w=3u
m:x8:18 n007 x8:nand 0 0 x8:nfet l=0.6u w=1.5u
m:x9:1 vdd x9:na x9:n001 vdd x9:pfet l=0.6u w=6u
m:x9:2 x9:n001 b9 p9 vdd x9:pfet l=0.6u w=6u
m:x9:3 vdd a9 x9:n002 vdd x9:pfet l=0.6u w=6u
m:x9:4 x9:n002 x9:nb p9 vdd x9:pfet l=0.6u w=6u
m:x9:5 p9 b9 x9:n004 0 x9:nfet l=0.6u w=3u
m:x9:6 x9:n004 a9 0 0 x9:nfet l=0.6u w=3u
m:x9:7 p9 x9:nb x9:n005 0 x9:nfet l=0.6u w=3u
m:x9:8 x9:n005 x9:na 0 0 x9:nfet l=0.6u w=3u
m:x9:9 vdd b9 x9:nb vdd x9:pfet l=0.6u w=3u
m:x9:10 x9:nb b9 0 0 x9:nfet l=0.6u w=1.5u
m:x9:11 vdd a9 x9:na vdd x9:pfet l=0.6u w=3u
m:x9:12 x9:na a9 0 0 x9:nfet l=0.6u w=1.5u
m:x9:13 x9:nand b9 x9:n003 0 x9:nfet l=0.6u w=3u
m:x9:14 x9:n003 a9 0 0 x9:nfet l=0.6u w=3u
m:x9:15 vdd a9 x9:nand vdd x9:pfet l=0.6u w=3u
m:x9:16 vdd b9 x9:nand vdd x9:pfet l=0.6u w=3u
m:x9:17 vdd x9:nand n006 vdd x9:pfet l=0.6u w=3u
m:x9:18 n006 x9:nand 0 0 x9:nfet l=0.6u w=1.5u
m:x10:1 vdd x10:na x10:n001 vdd x10:pfet l=0.6u w=6u
m:x10:2 x10:n001 b10 p10 vdd x10:pfet l=0.6u w=6u
m:x10:3 vdd a10 x10:n002 vdd x10:pfet l=0.6u w=6u
m:x10:4 x10:n002 x10:nb p10 vdd x10:pfet l=0.6u w=6u
m:x10:5 p10 b10 x10:n004 0 x10:nfet l=0.6u w=3u
m:x10:6 x10:n004 a10 0 0 x10:nfet l=0.6u w=3u
m:x10:7 p10 x10:nb x10:n005 0 x10:nfet l=0.6u w=3u
m:x10:8 x10:n005 x10:na 0 0 x10:nfet l=0.6u w=3u
m:x10:9 vdd b10 x10:nb vdd x10:pfet l=0.6u w=3u
m:x10:10 x10:nb b10 0 0 x10:nfet l=0.6u w=1.5u
m:x10:11 vdd a10 x10:na vdd x10:pfet l=0.6u w=3u
m:x10:12 x10:na a10 0 0 x10:nfet l=0.6u w=1.5u
m:x10:13 x10:nand b10 x10:n003 0 x10:nfet l=0.6u w=3u
m:x10:14 x10:n003 a10 0 0 x10:nfet l=0.6u w=3u
m:x10:15 vdd a10 x10:nand vdd x10:pfet l=0.6u w=3u
m:x10:16 vdd b10 x10:nand vdd x10:pfet l=0.6u w=3u
m:x10:17 vdd x10:nand n005 vdd x10:pfet l=0.6u w=3u
m:x10:18 n005 x10:nand 0 0 x10:nfet l=0.6u w=1.5u
m:x11:1 vdd x11:na x11:n001 vdd x11:pfet l=0.6u w=6u
m:x11:2 x11:n001 b11 p11 vdd x11:pfet l=0.6u w=6u
m:x11:3 vdd a11 x11:n002 vdd x11:pfet l=0.6u w=6u
m:x11:4 x11:n002 x11:nb p11 vdd x11:pfet l=0.6u w=6u
m:x11:5 p11 b11 x11:n004 0 x11:nfet l=0.6u w=3u
m:x11:6 x11:n004 a11 0 0 x11:nfet l=0.6u w=3u
m:x11:7 p11 x11:nb x11:n005 0 x11:nfet l=0.6u w=3u
m:x11:8 x11:n005 x11:na 0 0 x11:nfet l=0.6u w=3u
m:x11:9 vdd b11 x11:nb vdd x11:pfet l=0.6u w=3u
m:x11:10 x11:nb b11 0 0 x11:nfet l=0.6u w=1.5u
m:x11:11 vdd a11 x11:na vdd x11:pfet l=0.6u w=3u
m:x11:12 x11:na a11 0 0 x11:nfet l=0.6u w=1.5u
m:x11:13 x11:nand b11 x11:n003 0 x11:nfet l=0.6u w=3u
m:x11:14 x11:n003 a11 0 0 x11:nfet l=0.6u w=3u
m:x11:15 vdd a11 x11:nand vdd x11:pfet l=0.6u w=3u
m:x11:16 vdd b11 x11:nand vdd x11:pfet l=0.6u w=3u
m:x11:17 vdd x11:nand n004 vdd x11:pfet l=0.6u w=3u
m:x11:18 n004 x11:nand 0 0 x11:nfet l=0.6u w=1.5u
m:x12:1 vdd x12:na x12:n001 vdd x12:pfet l=0.6u w=6u
m:x12:2 x12:n001 b12 p12 vdd x12:pfet l=0.6u w=6u
m:x12:3 vdd a12 x12:n002 vdd x12:pfet l=0.6u w=6u
m:x12:4 x12:n002 x12:nb p12 vdd x12:pfet l=0.6u w=6u
m:x12:5 p12 b12 x12:n004 0 x12:nfet l=0.6u w=3u
m:x12:6 x12:n004 a12 0 0 x12:nfet l=0.6u w=3u
m:x12:7 p12 x12:nb x12:n005 0 x12:nfet l=0.6u w=3u
m:x12:8 x12:n005 x12:na 0 0 x12:nfet l=0.6u w=3u
m:x12:9 vdd b12 x12:nb vdd x12:pfet l=0.6u w=3u
m:x12:10 x12:nb b12 0 0 x12:nfet l=0.6u w=1.5u
m:x12:11 vdd a12 x12:na vdd x12:pfet l=0.6u w=3u
m:x12:12 x12:na a12 0 0 x12:nfet l=0.6u w=1.5u
m:x12:13 x12:nand b12 x12:n003 0 x12:nfet l=0.6u w=3u
m:x12:14 x12:n003 a12 0 0 x12:nfet l=0.6u w=3u
m:x12:15 vdd a12 x12:nand vdd x12:pfet l=0.6u w=3u
m:x12:16 vdd b12 x12:nand vdd x12:pfet l=0.6u w=3u
m:x12:17 vdd x12:nand n003 vdd x12:pfet l=0.6u w=3u
m:x12:18 n003 x12:nand 0 0 x12:nfet l=0.6u w=1.5u
m:x13:1 vdd x13:na x13:n001 vdd x13:pfet l=0.6u w=6u
m:x13:2 x13:n001 b13 p13 vdd x13:pfet l=0.6u w=6u
m:x13:3 vdd a13 x13:n002 vdd x13:pfet l=0.6u w=6u
m:x13:4 x13:n002 x13:nb p13 vdd x13:pfet l=0.6u w=6u
m:x13:5 p13 b13 x13:n004 0 x13:nfet l=0.6u w=3u
m:x13:6 x13:n004 a13 0 0 x13:nfet l=0.6u w=3u
m:x13:7 p13 x13:nb x13:n005 0 x13:nfet l=0.6u w=3u
m:x13:8 x13:n005 x13:na 0 0 x13:nfet l=0.6u w=3u
m:x13:9 vdd b13 x13:nb vdd x13:pfet l=0.6u w=3u
m:x13:10 x13:nb b13 0 0 x13:nfet l=0.6u w=1.5u
m:x13:11 vdd a13 x13:na vdd x13:pfet l=0.6u w=3u
m:x13:12 x13:na a13 0 0 x13:nfet l=0.6u w=1.5u
m:x13:13 x13:nand b13 x13:n003 0 x13:nfet l=0.6u w=3u
m:x13:14 x13:n003 a13 0 0 x13:nfet l=0.6u w=3u
m:x13:15 vdd a13 x13:nand vdd x13:pfet l=0.6u w=3u
m:x13:16 vdd b13 x13:nand vdd x13:pfet l=0.6u w=3u
m:x13:17 vdd x13:nand n002 vdd x13:pfet l=0.6u w=3u
m:x13:18 n002 x13:nand 0 0 x13:nfet l=0.6u w=1.5u
m:x14:1 vdd x14:na x14:n001 vdd x14:pfet l=0.6u w=6u
m:x14:2 x14:n001 b14 p14 vdd x14:pfet l=0.6u w=6u
m:x14:3 vdd a14 x14:n002 vdd x14:pfet l=0.6u w=6u
m:x14:4 x14:n002 x14:nb p14 vdd x14:pfet l=0.6u w=6u
m:x14:5 p14 b14 x14:n004 0 x14:nfet l=0.6u w=3u
m:x14:6 x14:n004 a14 0 0 x14:nfet l=0.6u w=3u
m:x14:7 p14 x14:nb x14:n005 0 x14:nfet l=0.6u w=3u
m:x14:8 x14:n005 x14:na 0 0 x14:nfet l=0.6u w=3u
m:x14:9 vdd b14 x14:nb vdd x14:pfet l=0.6u w=3u
m:x14:10 x14:nb b14 0 0 x14:nfet l=0.6u w=1.5u
m:x14:11 vdd a14 x14:na vdd x14:pfet l=0.6u w=3u
m:x14:12 x14:na a14 0 0 x14:nfet l=0.6u w=1.5u
m:x14:13 x14:nand b14 x14:n003 0 x14:nfet l=0.6u w=3u
m:x14:14 x14:n003 a14 0 0 x14:nfet l=0.6u w=3u
m:x14:15 vdd a14 x14:nand vdd x14:pfet l=0.6u w=3u
m:x14:16 vdd b14 x14:nand vdd x14:pfet l=0.6u w=3u
m:x14:17 vdd x14:nand n001 vdd x14:pfet l=0.6u w=3u
m:x14:18 n001 x14:nand 0 0 x14:nfet l=0.6u w=1.5u
m:x15:1 vdd x15:na x15:n001 vdd x15:pfet l=0.6u w=6u
m:x15:2 x15:n001 b15 p15 vdd x15:pfet l=0.6u w=6u
m:x15:3 vdd a15 x15:n002 vdd x15:pfet l=0.6u w=6u
m:x15:4 x15:n002 x15:nb p15 vdd x15:pfet l=0.6u w=6u
m:x15:5 p15 b15 x15:n004 0 x15:nfet l=0.6u w=3u
m:x15:6 x15:n004 a15 0 0 x15:nfet l=0.6u w=3u
m:x15:7 p15 x15:nb x15:n005 0 x15:nfet l=0.6u w=3u
m:x15:8 x15:n005 x15:na 0 0 x15:nfet l=0.6u w=3u
m:x15:9 vdd b15 x15:nb vdd x15:pfet l=0.6u w=3u
m:x15:10 x15:nb b15 0 0 x15:nfet l=0.6u w=1.5u
m:x15:11 vdd a15 x15:na vdd x15:pfet l=0.6u w=3u
m:x15:12 x15:na a15 0 0 x15:nfet l=0.6u w=1.5u
m:x15:13 x15:nand b15 x15:n003 0 x15:nfet l=0.6u w=3u
m:x15:14 x15:n003 a15 0 0 x15:nfet l=0.6u w=3u
m:x15:15 vdd a15 x15:nand vdd x15:pfet l=0.6u w=3u
m:x15:16 vdd b15 x15:nand vdd x15:pfet l=0.6u w=3u
m:x15:17 vdd x15:nand n015 vdd x15:pfet l=0.6u w=3u
m:x15:18 n015 x15:nand 0 0 x15:nfet l=0.6u w=1.5u
m:x17:1 vdd x17:n001 n039 vdd x17:pfet l=0.6u w=3u
m:x17:2 n039 x17:n001 0 0 x17:nfet l=0.6u w=1.5u
m:x17:3 vdd cin x17:n001 vdd x17:pfet l=0.6u w=3u
m:x17:4 x17:n001 cin 0 0 x17:nfet l=0.6u w=1.5u
m:x18:1 vdd p1 x18:nb vdd x18:pfet l=0.6u w=3u
m:x18:2 x18:nb p1 0 0 x18:nfet l=0.6u w=1.5u
m:x18:3 vdd cin x18:na vdd x18:pfet l=0.6u w=3u
m:x18:4 x18:na cin 0 0 x18:nfet l=0.6u w=1.5u
m:x18:5 vdd n014 x18:nc vdd x18:pfet l=0.6u w=3u
m:x18:6 x18:nc n014 0 0 x18:nfet l=0.6u w=1.5u
m:x18:7 vdd x18:nc n036 vdd x18:pfet l=0.6u w=3u
m:x18:8 vdd x18:na x18:n001 vdd x18:pfet l=0.6u w=3u
m:x18:9 x18:n001 x18:nb n036 vdd x18:pfet l=0.6u w=3u
m:x18:10 n036 x18:na x18:n002 0 x18:nfet l=0.6u w=1.5u
m:x18:11 n036 x18:nb x18:n002 0 x18:nfet l=0.6u w=1.5u
m:x18:12 x18:n002 x18:nc 0 0 x18:nfet l=0.6u w=1.5u
m:x19:1 vdd p2 x19:nb vdd x19:pfet l=0.6u w=3u
m:x19:2 x19:nb p2 0 0 x19:nfet l=0.6u w=1.5u
m:x19:3 vdd n014 x19:na vdd x19:pfet l=0.6u w=3u
m:x19:4 x19:na n014 0 0 x19:nfet l=0.6u w=1.5u
m:x19:5 vdd n013 x19:nc vdd x19:pfet l=0.6u w=3u
m:x19:6 x19:nc n013 0 0 x19:nfet l=0.6u w=1.5u
m:x19:7 vdd x19:nc n030 vdd x19:pfet l=0.6u w=6u
m:x19:8 vdd x19:nb x19:n001 vdd x19:pfet l=0.6u w=6u
m:x19:9 x19:n001 x19:na n030 vdd x19:pfet l=0.6u w=6u
m:x19:10 n030 x19:na x19:n004 0 x19:nfet l=0.6u w=3u
m:x19:11 n030 x19:nb x19:n004 0 x19:nfet l=0.6u w=3u
m:x19:12 x19:n004 x19:nc 0 0 x19:nfet l=0.6u w=3u
m:x19:13 x19:n003 p2 0 0 x19:nfet l=0.6u w=3u
m:x19:14 x19:n002 p1 x19:n003 0 x19:nfet l=0.6u w=3u
m:x19:15 vdd p2 x19:n002 vdd x19:pfet l=0.6u w=3u
m:x19:16 vdd p1 x19:n002 vdd x19:pfet l=0.6u w=3u
m:x19:17 vdd x19:n002 n033 vdd x19:pfet l=0.6u w=3u
m:x19:18 n033 x19:n002 0 0 x19:nfet l=0.6u w=1.5u
m:x20:1 vdd p3 x20:nb vdd x20:pfet l=0.6u w=3u
m:x20:2 x20:nb p3 0 0 x20:nfet l=0.6u w=1.5u
m:x20:3 vdd n013 x20:na vdd x20:pfet l=0.6u w=3u
m:x20:4 x20:na n013 0 0 x20:nfet l=0.6u w=1.5u
m:x20:5 vdd n012 x20:nc vdd x20:pfet l=0.6u w=3u
m:x20:6 x20:nc n012 0 0 x20:nfet l=0.6u w=1.5u
m:x20:7 vdd x20:nc n024 vdd x20:pfet l=0.6u w=6u
m:x20:8 vdd x20:nb x20:n001 vdd x20:pfet l=0.6u w=6u
m:x20:9 x20:n001 x20:na n024 vdd x20:pfet l=0.6u w=6u
m:x20:10 n024 x20:na x20:n004 0 x20:nfet l=0.6u w=3u
m:x20:11 n024 x20:nb x20:n004 0 x20:nfet l=0.6u w=3u
m:x20:12 x20:n004 x20:nc 0 0 x20:nfet l=0.6u w=3u
m:x20:13 x20:n003 p3 0 0 x20:nfet l=0.6u w=3u
m:x20:14 x20:n002 p2 x20:n003 0 x20:nfet l=0.6u w=3u
m:x20:15 vdd p3 x20:n002 vdd x20:pfet l=0.6u w=3u
m:x20:16 vdd p2 x20:n002 vdd x20:pfet l=0.6u w=3u
m:x20:17 vdd x20:n002 n027 vdd x20:pfet l=0.6u w=3u
m:x20:18 n027 x20:n002 0 0 x20:nfet l=0.6u w=1.5u
m:x21:1 vdd p4 x21:nb vdd x21:pfet l=0.6u w=3u
m:x21:2 x21:nb p4 0 0 x21:nfet l=0.6u w=1.5u
m:x21:3 vdd n012 x21:na vdd x21:pfet l=0.6u w=3u
m:x21:4 x21:na n012 0 0 x21:nfet l=0.6u w=1.5u
m:x21:5 vdd n011 x21:nc vdd x21:pfet l=0.6u w=3u
m:x21:6 x21:nc n011 0 0 x21:nfet l=0.6u w=1.5u
m:x21:7 vdd x21:nc n018 vdd x21:pfet l=0.6u w=6u
m:x21:8 vdd x21:nb x21:n001 vdd x21:pfet l=0.6u w=6u
m:x21:9 x21:n001 x21:na n018 vdd x21:pfet l=0.6u w=6u
m:x21:10 n018 x21:na x21:n004 0 x21:nfet l=0.6u w=3u
m:x21:11 n018 x21:nb x21:n004 0 x21:nfet l=0.6u w=3u
m:x21:12 x21:n004 x21:nc 0 0 x21:nfet l=0.6u w=3u
m:x21:13 x21:n003 p4 0 0 x21:nfet l=0.6u w=3u
m:x21:14 x21:n002 p3 x21:n003 0 x21:nfet l=0.6u w=3u
m:x21:15 vdd p4 x21:n002 vdd x21:pfet l=0.6u w=3u
m:x21:16 vdd p3 x21:n002 vdd x21:pfet l=0.6u w=3u
m:x21:17 vdd x21:n002 n021 vdd x21:pfet l=0.6u w=3u
m:x21:18 n021 x21:n002 0 0 x21:nfet l=0.6u w=1.5u
m:x22:1 vdd p5 x22:nb vdd x22:pfet l=0.6u w=3u
m:x22:2 x22:nb p5 0 0 x22:nfet l=0.6u w=1.5u
m:x22:3 vdd n011 x22:na vdd x22:pfet l=0.6u w=3u
m:x22:4 x22:na n011 0 0 x22:nfet l=0.6u w=1.5u
m:x22:5 vdd n010 x22:nc vdd x22:pfet l=0.6u w=3u
m:x22:6 x22:nc n010 0 0 x22:nfet l=0.6u w=1.5u
m:x22:7 vdd x22:nc n035 vdd x22:pfet l=0.6u w=6u
m:x22:8 vdd x22:nb x22:n001 vdd x22:pfet l=0.6u w=6u
m:x22:9 x22:n001 x22:na n035 vdd x22:pfet l=0.6u w=6u
m:x22:10 n035 x22:na x22:n004 0 x22:nfet l=0.6u w=3u
m:x22:11 n035 x22:nb x22:n004 0 x22:nfet l=0.6u w=3u
m:x22:12 x22:n004 x22:nc 0 0 x22:nfet l=0.6u w=3u
m:x22:13 x22:n003 p5 0 0 x22:nfet l=0.6u w=3u
m:x22:14 x22:n002 p4 x22:n003 0 x22:nfet l=0.6u w=3u
m:x22:15 vdd p5 x22:n002 vdd x22:pfet l=0.6u w=3u
m:x22:16 vdd p4 x22:n002 vdd x22:pfet l=0.6u w=3u
m:x22:17 vdd x22:n002 n038 vdd x22:pfet l=0.6u w=3u
m:x22:18 n038 x22:n002 0 0 x22:nfet l=0.6u w=1.5u
m:x23:1 vdd p6 x23:nb vdd x23:pfet l=0.6u w=3u
m:x23:2 x23:nb p6 0 0 x23:nfet l=0.6u w=1.5u
m:x23:3 vdd n010 x23:na vdd x23:pfet l=0.6u w=3u
m:x23:4 x23:na n010 0 0 x23:nfet l=0.6u w=1.5u
m:x23:5 vdd n009 x23:nc vdd x23:pfet l=0.6u w=3u
m:x23:6 x23:nc n009 0 0 x23:nfet l=0.6u w=1.5u
m:x23:7 vdd x23:nc n029 vdd x23:pfet l=0.6u w=6u
m:x23:8 vdd x23:nb x23:n001 vdd x23:pfet l=0.6u w=6u
m:x23:9 x23:n001 x23:na n029 vdd x23:pfet l=0.6u w=6u
m:x23:10 n029 x23:na x23:n004 0 x23:nfet l=0.6u w=3u
m:x23:11 n029 x23:nb x23:n004 0 x23:nfet l=0.6u w=3u
m:x23:12 x23:n004 x23:nc 0 0 x23:nfet l=0.6u w=3u
m:x23:13 x23:n003 p6 0 0 x23:nfet l=0.6u w=3u
m:x23:14 x23:n002 p5 x23:n003 0 x23:nfet l=0.6u w=3u
m:x23:15 vdd p6 x23:n002 vdd x23:pfet l=0.6u w=3u
m:x23:16 vdd p5 x23:n002 vdd x23:pfet l=0.6u w=3u
m:x23:17 vdd x23:n002 n032 vdd x23:pfet l=0.6u w=3u
m:x23:18 n032 x23:n002 0 0 x23:nfet l=0.6u w=1.5u
m:x24:1 vdd p7 x24:nb vdd x24:pfet l=0.6u w=3u
m:x24:2 x24:nb p7 0 0 x24:nfet l=0.6u w=1.5u
m:x24:3 vdd n009 x24:na vdd x24:pfet l=0.6u w=3u
m:x24:4 x24:na n009 0 0 x24:nfet l=0.6u w=1.5u
m:x24:5 vdd n008 x24:nc vdd x24:pfet l=0.6u w=3u
m:x24:6 x24:nc n008 0 0 x24:nfet l=0.6u w=1.5u
m:x24:7 vdd x24:nc n023 vdd x24:pfet l=0.6u w=6u
m:x24:8 vdd x24:nb x24:n001 vdd x24:pfet l=0.6u w=6u
m:x24:9 x24:n001 x24:na n023 vdd x24:pfet l=0.6u w=6u
m:x24:10 n023 x24:na x24:n004 0 x24:nfet l=0.6u w=3u
m:x24:11 n023 x24:nb x24:n004 0 x24:nfet l=0.6u w=3u
m:x24:12 x24:n004 x24:nc 0 0 x24:nfet l=0.6u w=3u
m:x24:13 x24:n003 p7 0 0 x24:nfet l=0.6u w=3u
m:x24:14 x24:n002 p6 x24:n003 0 x24:nfet l=0.6u w=3u
m:x24:15 vdd p7 x24:n002 vdd x24:pfet l=0.6u w=3u
m:x24:16 vdd p6 x24:n002 vdd x24:pfet l=0.6u w=3u
m:x24:17 vdd x24:n002 n026 vdd x24:pfet l=0.6u w=3u
m:x24:18 n026 x24:n002 0 0 x24:nfet l=0.6u w=1.5u
m:x25:1 vdd p8 x25:nb vdd x25:pfet l=0.6u w=3u
m:x25:2 x25:nb p8 0 0 x25:nfet l=0.6u w=1.5u
m:x25:3 vdd n008 x25:na vdd x25:pfet l=0.6u w=3u
m:x25:4 x25:na n008 0 0 x25:nfet l=0.6u w=1.5u
m:x25:5 vdd n007 x25:nc vdd x25:pfet l=0.6u w=3u
m:x25:6 x25:nc n007 0 0 x25:nfet l=0.6u w=1.5u
m:x25:7 vdd x25:nc n017 vdd x25:pfet l=0.6u w=6u
m:x25:8 vdd x25:nb x25:n001 vdd x25:pfet l=0.6u w=6u
m:x25:9 x25:n001 x25:na n017 vdd x25:pfet l=0.6u w=6u
m:x25:10 n017 x25:na x25:n004 0 x25:nfet l=0.6u w=3u
m:x25:11 n017 x25:nb x25:n004 0 x25:nfet l=0.6u w=3u
m:x25:12 x25:n004 x25:nc 0 0 x25:nfet l=0.6u w=3u
m:x25:13 x25:n003 p8 0 0 x25:nfet l=0.6u w=3u
m:x25:14 x25:n002 p7 x25:n003 0 x25:nfet l=0.6u w=3u
m:x25:15 vdd p8 x25:n002 vdd x25:pfet l=0.6u w=3u
m:x25:16 vdd p7 x25:n002 vdd x25:pfet l=0.6u w=3u
m:x25:17 vdd x25:n002 n020 vdd x25:pfet l=0.6u w=3u
m:x25:18 n020 x25:n002 0 0 x25:nfet l=0.6u w=1.5u
m:x26:1 vdd p9 x26:nb vdd x26:pfet l=0.6u w=3u
m:x26:2 x26:nb p9 0 0 x26:nfet l=0.6u w=1.5u
m:x26:3 vdd n007 x26:na vdd x26:pfet l=0.6u w=3u
m:x26:4 x26:na n007 0 0 x26:nfet l=0.6u w=1.5u
m:x26:5 vdd n006 x26:nc vdd x26:pfet l=0.6u w=3u
m:x26:6 x26:nc n006 0 0 x26:nfet l=0.6u w=1.5u
m:x26:7 vdd x26:nc n034 vdd x26:pfet l=0.6u w=6u
m:x26:8 vdd x26:nb x26:n001 vdd x26:pfet l=0.6u w=6u
m:x26:9 x26:n001 x26:na n034 vdd x26:pfet l=0.6u w=6u
m:x26:10 n034 x26:na x26:n004 0 x26:nfet l=0.6u w=3u
m:x26:11 n034 x26:nb x26:n004 0 x26:nfet l=0.6u w=3u
m:x26:12 x26:n004 x26:nc 0 0 x26:nfet l=0.6u w=3u
m:x26:13 x26:n003 p9 0 0 x26:nfet l=0.6u w=3u
m:x26:14 x26:n002 p8 x26:n003 0 x26:nfet l=0.6u w=3u
m:x26:15 vdd p9 x26:n002 vdd x26:pfet l=0.6u w=3u
m:x26:16 vdd p8 x26:n002 vdd x26:pfet l=0.6u w=3u
m:x26:17 vdd x26:n002 n037 vdd x26:pfet l=0.6u w=3u
m:x26:18 n037 x26:n002 0 0 x26:nfet l=0.6u w=1.5u
m:x27:1 vdd p10 x27:nb vdd x27:pfet l=0.6u w=3u
m:x27:2 x27:nb p10 0 0 x27:nfet l=0.6u w=1.5u
m:x27:3 vdd n006 x27:na vdd x27:pfet l=0.6u w=3u
m:x27:4 x27:na n006 0 0 x27:nfet l=0.6u w=1.5u
m:x27:5 vdd n005 x27:nc vdd x27:pfet l=0.6u w=3u
m:x27:6 x27:nc n005 0 0 x27:nfet l=0.6u w=1.5u
m:x27:7 vdd x27:nc n028 vdd x27:pfet l=0.6u w=6u
m:x27:8 vdd x27:nb x27:n001 vdd x27:pfet l=0.6u w=6u
m:x27:9 x27:n001 x27:na n028 vdd x27:pfet l=0.6u w=6u
m:x27:10 n028 x27:na x27:n004 0 x27:nfet l=0.6u w=3u
m:x27:11 n028 x27:nb x27:n004 0 x27:nfet l=0.6u w=3u
m:x27:12 x27:n004 x27:nc 0 0 x27:nfet l=0.6u w=3u
m:x27:13 x27:n003 p10 0 0 x27:nfet l=0.6u w=3u
m:x27:14 x27:n002 p9 x27:n003 0 x27:nfet l=0.6u w=3u
m:x27:15 vdd p10 x27:n002 vdd x27:pfet l=0.6u w=3u
m:x27:16 vdd p9 x27:n002 vdd x27:pfet l=0.6u w=3u
m:x27:17 vdd x27:n002 n031 vdd x27:pfet l=0.6u w=3u
m:x27:18 n031 x27:n002 0 0 x27:nfet l=0.6u w=1.5u
m:x28:1 vdd p11 x28:nb vdd x28:pfet l=0.6u w=3u
m:x28:2 x28:nb p11 0 0 x28:nfet l=0.6u w=1.5u
m:x28:3 vdd n005 x28:na vdd x28:pfet l=0.6u w=3u
m:x28:4 x28:na n005 0 0 x28:nfet l=0.6u w=1.5u
m:x28:5 vdd n004 x28:nc vdd x28:pfet l=0.6u w=3u
m:x28:6 x28:nc n004 0 0 x28:nfet l=0.6u w=1.5u
m:x28:7 vdd x28:nc n022 vdd x28:pfet l=0.6u w=6u
m:x28:8 vdd x28:nb x28:n001 vdd x28:pfet l=0.6u w=6u
m:x28:9 x28:n001 x28:na n022 vdd x28:pfet l=0.6u w=6u
m:x28:10 n022 x28:na x28:n004 0 x28:nfet l=0.6u w=3u
m:x28:11 n022 x28:nb x28:n004 0 x28:nfet l=0.6u w=3u
m:x28:12 x28:n004 x28:nc 0 0 x28:nfet l=0.6u w=3u
m:x28:13 x28:n003 p11 0 0 x28:nfet l=0.6u w=3u
m:x28:14 x28:n002 p10 x28:n003 0 x28:nfet l=0.6u w=3u
m:x28:15 vdd p11 x28:n002 vdd x28:pfet l=0.6u w=3u
m:x28:16 vdd p10 x28:n002 vdd x28:pfet l=0.6u w=3u
m:x28:17 vdd x28:n002 n025 vdd x28:pfet l=0.6u w=3u
m:x28:18 n025 x28:n002 0 0 x28:nfet l=0.6u w=1.5u
m:x29:1 vdd p12 x29:nb vdd x29:pfet l=0.6u w=3u
m:x29:2 x29:nb p12 0 0 x29:nfet l=0.6u w=1.5u
m:x29:3 vdd n004 x29:na vdd x29:pfet l=0.6u w=3u
m:x29:4 x29:na n004 0 0 x29:nfet l=0.6u w=1.5u
m:x29:5 vdd n003 x29:nc vdd x29:pfet l=0.6u w=3u
m:x29:6 x29:nc n003 0 0 x29:nfet l=0.6u w=1.5u
m:x29:7 vdd x29:nc n016 vdd x29:pfet l=0.6u w=6u
m:x29:8 vdd x29:nb x29:n001 vdd x29:pfet l=0.6u w=6u
m:x29:9 x29:n001 x29:na n016 vdd x29:pfet l=0.6u w=6u
m:x29:10 n016 x29:na x29:n004 0 x29:nfet l=0.6u w=3u
m:x29:11 n016 x29:nb x29:n004 0 x29:nfet l=0.6u w=3u
m:x29:12 x29:n004 x29:nc 0 0 x29:nfet l=0.6u w=3u
m:x29:13 x29:n003 p12 0 0 x29:nfet l=0.6u w=3u
m:x29:14 x29:n002 p11 x29:n003 0 x29:nfet l=0.6u w=3u
m:x29:15 vdd p12 x29:n002 vdd x29:pfet l=0.6u w=3u
m:x29:16 vdd p11 x29:n002 vdd x29:pfet l=0.6u w=3u
m:x29:17 vdd x29:n002 n019 vdd x29:pfet l=0.6u w=3u
m:x29:18 n019 x29:n002 0 0 x29:nfet l=0.6u w=1.5u
m:x30:1 vdd p13 x30:nb vdd x30:pfet l=0.6u w=3u
m:x30:2 x30:nb p13 0 0 x30:nfet l=0.6u w=1.5u
m:x30:3 vdd n003 x30:na vdd x30:pfet l=0.6u w=3u
m:x30:4 x30:na n003 0 0 x30:nfet l=0.6u w=1.5u
m:x30:5 vdd n002 x30:nc vdd x30:pfet l=0.6u w=3u
m:x30:6 x30:nc n002 0 0 x30:nfet l=0.6u w=1.5u
m:x30:7 vdd x30:nc n044 vdd x30:pfet l=0.6u w=6u
m:x30:8 vdd x30:nb x30:n001 vdd x30:pfet l=0.6u w=6u
m:x30:9 x30:n001 x30:na n044 vdd x30:pfet l=0.6u w=6u
m:x30:10 n044 x30:na x30:n004 0 x30:nfet l=0.6u w=3u
m:x30:11 n044 x30:nb x30:n004 0 x30:nfet l=0.6u w=3u
m:x30:12 x30:n004 x30:nc 0 0 x30:nfet l=0.6u w=3u
m:x30:13 x30:n003 p13 0 0 x30:nfet l=0.6u w=3u
m:x30:14 x30:n002 p12 x30:n003 0 x30:nfet l=0.6u w=3u
m:x30:15 vdd p13 x30:n002 vdd x30:pfet l=0.6u w=3u
m:x30:16 vdd p12 x30:n002 vdd x30:pfet l=0.6u w=3u
m:x30:17 vdd x30:n002 n045 vdd x30:pfet l=0.6u w=3u
m:x30:18 n045 x30:n002 0 0 x30:nfet l=0.6u w=1.5u
m:x31:1 vdd p14 x31:nb vdd x31:pfet l=0.6u w=3u
m:x31:2 x31:nb p14 0 0 x31:nfet l=0.6u w=1.5u
m:x31:3 vdd n002 x31:na vdd x31:pfet l=0.6u w=3u
m:x31:4 x31:na n002 0 0 x31:nfet l=0.6u w=1.5u
m:x31:5 vdd n001 x31:nc vdd x31:pfet l=0.6u w=3u
m:x31:6 x31:nc n001 0 0 x31:nfet l=0.6u w=1.5u
m:x31:7 vdd x31:nc n042 vdd x31:pfet l=0.6u w=6u
m:x31:8 vdd x31:nb x31:n001 vdd x31:pfet l=0.6u w=6u
m:x31:9 x31:n001 x31:na n042 vdd x31:pfet l=0.6u w=6u
m:x31:10 n042 x31:na x31:n004 0 x31:nfet l=0.6u w=3u
m:x31:11 n042 x31:nb x31:n004 0 x31:nfet l=0.6u w=3u
m:x31:12 x31:n004 x31:nc 0 0 x31:nfet l=0.6u w=3u
m:x31:13 x31:n003 p14 0 0 x31:nfet l=0.6u w=3u
m:x31:14 x31:n002 p13 x31:n003 0 x31:nfet l=0.6u w=3u
m:x31:15 vdd p14 x31:n002 vdd x31:pfet l=0.6u w=3u
m:x31:16 vdd p13 x31:n002 vdd x31:pfet l=0.6u w=3u
m:x31:17 vdd x31:n002 n043 vdd x31:pfet l=0.6u w=3u
m:x31:18 n043 x31:n002 0 0 x31:nfet l=0.6u w=1.5u
m:x34:1 vdd x34:n001 n060 vdd x34:pfet l=0.6u w=3u
m:x34:2 n060 x34:n001 0 0 x34:nfet l=0.6u w=1.5u
m:x34:3 vdd n036 x34:n001 vdd x34:pfet l=0.6u w=3u
m:x34:4 x34:n001 n036 0 0 x34:nfet l=0.6u w=1.5u
m:x35:1 vdd n033 x35:nb vdd x35:pfet l=0.6u w=3u
m:x35:2 x35:nb n033 0 0 x35:nfet l=0.6u w=1.5u
m:x35:3 vdd n039 x35:na vdd x35:pfet l=0.6u w=3u
m:x35:4 x35:na n039 0 0 x35:nfet l=0.6u w=1.5u
m:x35:5 vdd n030 x35:nc vdd x35:pfet l=0.6u w=3u
m:x35:6 x35:nc n030 0 0 x35:nfet l=0.6u w=1.5u
m:x35:7 vdd x35:nc n057 vdd x35:pfet l=0.6u w=3u
m:x35:8 vdd x35:na x35:n001 vdd x35:pfet l=0.6u w=3u
m:x35:9 x35:n001 x35:nb n057 vdd x35:pfet l=0.6u w=3u
m:x35:10 n057 x35:na x35:n002 0 x35:nfet l=0.6u w=1.5u
m:x35:11 n057 x35:nb x35:n002 0 x35:nfet l=0.6u w=1.5u
m:x35:12 x35:n002 x35:nc 0 0 x35:nfet l=0.6u w=1.5u
m:x36:1 vdd n027 x36:nb vdd x36:pfet l=0.6u w=3u
m:x36:2 x36:nb n027 0 0 x36:nfet l=0.6u w=1.5u
m:x36:3 vdd n036 x36:na vdd x36:pfet l=0.6u w=3u
m:x36:4 x36:na n036 0 0 x36:nfet l=0.6u w=1.5u
m:x36:5 vdd n024 x36:nc vdd x36:pfet l=0.6u w=3u
m:x36:6 x36:nc n024 0 0 x36:nfet l=0.6u w=1.5u
m:x36:7 vdd x36:nc n054 vdd x36:pfet l=0.6u w=3u
m:x36:8 vdd x36:na x36:n001 vdd x36:pfet l=0.6u w=3u
m:x36:9 x36:n001 x36:nb n054 vdd x36:pfet l=0.6u w=3u
m:x36:10 n054 x36:na x36:n002 0 x36:nfet l=0.6u w=1.5u
m:x36:11 n054 x36:nb x36:n002 0 x36:nfet l=0.6u w=1.5u
m:x36:12 x36:n002 x36:nc 0 0 x36:nfet l=0.6u w=1.5u
m:x37:1 vdd n021 x37:nb vdd x37:pfet l=0.6u w=3u
m:x37:2 x37:nb n021 0 0 x37:nfet l=0.6u w=1.5u
m:x37:3 vdd n030 x37:na vdd x37:pfet l=0.6u w=3u
m:x37:4 x37:na n030 0 0 x37:nfet l=0.6u w=1.5u
m:x37:5 vdd n018 x37:nc vdd x37:pfet l=0.6u w=3u
m:x37:6 x37:nc n018 0 0 x37:nfet l=0.6u w=1.5u
m:x37:7 vdd x37:nc n062 vdd x37:pfet l=0.6u w=6u
m:x37:8 vdd x37:nb x37:n001 vdd x37:pfet l=0.6u w=6u
m:x37:9 x37:n001 x37:na n062 vdd x37:pfet l=0.6u w=6u
m:x37:10 n062 x37:na x37:n004 0 x37:nfet l=0.6u w=3u
m:x37:11 n062 x37:nb x37:n004 0 x37:nfet l=0.6u w=3u
m:x37:12 x37:n004 x37:nc 0 0 x37:nfet l=0.6u w=3u
m:x37:13 x37:n003 n021 0 0 x37:nfet l=0.6u w=3u
m:x37:14 x37:n002 n033 x37:n003 0 x37:nfet l=0.6u w=3u
m:x37:15 vdd n021 x37:n002 vdd x37:pfet l=0.6u w=3u
m:x37:16 vdd n033 x37:n002 vdd x37:pfet l=0.6u w=3u
m:x37:17 vdd x37:n002 n064 vdd x37:pfet l=0.6u w=3u
m:x37:18 n064 x37:n002 0 0 x37:nfet l=0.6u w=1.5u
m:x38:1 vdd n038 x38:nb vdd x38:pfet l=0.6u w=3u
m:x38:2 x38:nb n038 0 0 x38:nfet l=0.6u w=1.5u
m:x38:3 vdd n024 x38:na vdd x38:pfet l=0.6u w=3u
m:x38:4 x38:na n024 0 0 x38:nfet l=0.6u w=1.5u
m:x38:5 vdd n035 x38:nc vdd x38:pfet l=0.6u w=3u
m:x38:6 x38:nc n035 0 0 x38:nfet l=0.6u w=1.5u
m:x38:7 vdd x38:nc n058 vdd x38:pfet l=0.6u w=6u
m:x38:8 vdd x38:nb x38:n001 vdd x38:pfet l=0.6u w=6u
m:x38:9 x38:n001 x38:na n058 vdd x38:pfet l=0.6u w=6u
m:x38:10 n058 x38:na x38:n004 0 x38:nfet l=0.6u w=3u
m:x38:11 n058 x38:nb x38:n004 0 x38:nfet l=0.6u w=3u
m:x38:12 x38:n004 x38:nc 0 0 x38:nfet l=0.6u w=3u
m:x38:13 x38:n003 n038 0 0 x38:nfet l=0.6u w=3u
m:x38:14 x38:n002 n027 x38:n003 0 x38:nfet l=0.6u w=3u
m:x38:15 vdd n038 x38:n002 vdd x38:pfet l=0.6u w=3u
m:x38:16 vdd n027 x38:n002 vdd x38:pfet l=0.6u w=3u
m:x38:17 vdd x38:n002 n059 vdd x38:pfet l=0.6u w=3u
m:x38:18 n059 x38:n002 0 0 x38:nfet l=0.6u w=1.5u
m:x39:1 vdd n032 x39:nb vdd x39:pfet l=0.6u w=3u
m:x39:2 x39:nb n032 0 0 x39:nfet l=0.6u w=1.5u
m:x39:3 vdd n018 x39:na vdd x39:pfet l=0.6u w=3u
m:x39:4 x39:na n018 0 0 x39:nfet l=0.6u w=1.5u
m:x39:5 vdd n029 x39:nc vdd x39:pfet l=0.6u w=3u
m:x39:6 x39:nc n029 0 0 x39:nfet l=0.6u w=1.5u
m:x39:7 vdd x39:nc n055 vdd x39:pfet l=0.6u w=6u
m:x39:8 vdd x39:nb x39:n001 vdd x39:pfet l=0.6u w=6u
m:x39:9 x39:n001 x39:na n055 vdd x39:pfet l=0.6u w=6u
m:x39:10 n055 x39:na x39:n004 0 x39:nfet l=0.6u w=3u
m:x39:11 n055 x39:nb x39:n004 0 x39:nfet l=0.6u w=3u
m:x39:12 x39:n004 x39:nc 0 0 x39:nfet l=0.6u w=3u
m:x39:13 x39:n003 n032 0 0 x39:nfet l=0.6u w=3u
m:x39:14 x39:n002 n021 x39:n003 0 x39:nfet l=0.6u w=3u
m:x39:15 vdd n032 x39:n002 vdd x39:pfet l=0.6u w=3u
m:x39:16 vdd n021 x39:n002 vdd x39:pfet l=0.6u w=3u
m:x39:17 vdd x39:n002 n056 vdd x39:pfet l=0.6u w=3u
m:x39:18 n056 x39:n002 0 0 x39:nfet l=0.6u w=1.5u
m:x40:1 vdd n026 x40:nb vdd x40:pfet l=0.6u w=3u
m:x40:2 x40:nb n026 0 0 x40:nfet l=0.6u w=1.5u
m:x40:3 vdd n035 x40:na vdd x40:pfet l=0.6u w=3u
m:x40:4 x40:na n035 0 0 x40:nfet l=0.6u w=1.5u
m:x40:5 vdd n023 x40:nc vdd x40:pfet l=0.6u w=3u
m:x40:6 x40:nc n023 0 0 x40:nfet l=0.6u w=1.5u
m:x40:7 vdd x40:nc n052 vdd x40:pfet l=0.6u w=6u
m:x40:8 vdd x40:nb x40:n001 vdd x40:pfet l=0.6u w=6u
m:x40:9 x40:n001 x40:na n052 vdd x40:pfet l=0.6u w=6u
m:x40:10 n052 x40:na x40:n004 0 x40:nfet l=0.6u w=3u
m:x40:11 n052 x40:nb x40:n004 0 x40:nfet l=0.6u w=3u
m:x40:12 x40:n004 x40:nc 0 0 x40:nfet l=0.6u w=3u
m:x40:13 x40:n003 n026 0 0 x40:nfet l=0.6u w=3u
m:x40:14 x40:n002 n038 x40:n003 0 x40:nfet l=0.6u w=3u
m:x40:15 vdd n026 x40:n002 vdd x40:pfet l=0.6u w=3u
m:x40:16 vdd n038 x40:n002 vdd x40:pfet l=0.6u w=3u
m:x40:17 vdd x40:n002 n053 vdd x40:pfet l=0.6u w=3u
m:x40:18 n053 x40:n002 0 0 x40:nfet l=0.6u w=1.5u
m:x41:1 vdd n020 x41:nb vdd x41:pfet l=0.6u w=3u
m:x41:2 x41:nb n020 0 0 x41:nfet l=0.6u w=1.5u
m:x41:3 vdd n029 x41:na vdd x41:pfet l=0.6u w=3u
m:x41:4 x41:na n029 0 0 x41:nfet l=0.6u w=1.5u
m:x41:5 vdd n017 x41:nc vdd x41:pfet l=0.6u w=3u
m:x41:6 x41:nc n017 0 0 x41:nfet l=0.6u w=1.5u
m:x41:7 vdd x41:nc n050 vdd x41:pfet l=0.6u w=6u
m:x41:8 vdd x41:nb x41:n001 vdd x41:pfet l=0.6u w=6u
m:x41:9 x41:n001 x41:na n050 vdd x41:pfet l=0.6u w=6u
m:x41:10 n050 x41:na x41:n004 0 x41:nfet l=0.6u w=3u
m:x41:11 n050 x41:nb x41:n004 0 x41:nfet l=0.6u w=3u
m:x41:12 x41:n004 x41:nc 0 0 x41:nfet l=0.6u w=3u
m:x41:13 x41:n003 n020 0 0 x41:nfet l=0.6u w=3u
m:x41:14 x41:n002 n032 x41:n003 0 x41:nfet l=0.6u w=3u
m:x41:15 vdd n020 x41:n002 vdd x41:pfet l=0.6u w=3u
m:x41:16 vdd n032 x41:n002 vdd x41:pfet l=0.6u w=3u
m:x41:17 vdd x41:n002 n051 vdd x41:pfet l=0.6u w=3u
m:x41:18 n051 x41:n002 0 0 x41:nfet l=0.6u w=1.5u
m:x42:1 vdd n037 x42:nb vdd x42:pfet l=0.6u w=3u
m:x42:2 x42:nb n037 0 0 x42:nfet l=0.6u w=1.5u
m:x42:3 vdd n023 x42:na vdd x42:pfet l=0.6u w=3u
m:x42:4 x42:na n023 0 0 x42:nfet l=0.6u w=1.5u
m:x42:5 vdd n034 x42:nc vdd x42:pfet l=0.6u w=3u
m:x42:6 x42:nc n034 0 0 x42:nfet l=0.6u w=1.5u
m:x42:7 vdd x42:nc n048 vdd x42:pfet l=0.6u w=6u
m:x42:8 vdd x42:nb x42:n001 vdd x42:pfet l=0.6u w=6u
m:x42:9 x42:n001 x42:na n048 vdd x42:pfet l=0.6u w=6u
m:x42:10 n048 x42:na x42:n004 0 x42:nfet l=0.6u w=3u
m:x42:11 n048 x42:nb x42:n004 0 x42:nfet l=0.6u w=3u
m:x42:12 x42:n004 x42:nc 0 0 x42:nfet l=0.6u w=3u
m:x42:13 x42:n003 n037 0 0 x42:nfet l=0.6u w=3u
m:x42:14 x42:n002 n026 x42:n003 0 x42:nfet l=0.6u w=3u
m:x42:15 vdd n037 x42:n002 vdd x42:pfet l=0.6u w=3u
m:x42:16 vdd n026 x42:n002 vdd x42:pfet l=0.6u w=3u
m:x42:17 vdd x42:n002 n049 vdd x42:pfet l=0.6u w=3u
m:x42:18 n049 x42:n002 0 0 x42:nfet l=0.6u w=1.5u
m:x43:1 vdd n031 x43:nb vdd x43:pfet l=0.6u w=3u
m:x43:2 x43:nb n031 0 0 x43:nfet l=0.6u w=1.5u
m:x43:3 vdd n017 x43:na vdd x43:pfet l=0.6u w=3u
m:x43:4 x43:na n017 0 0 x43:nfet l=0.6u w=1.5u
m:x43:5 vdd n028 x43:nc vdd x43:pfet l=0.6u w=3u
m:x43:6 x43:nc n028 0 0 x43:nfet l=0.6u w=1.5u
m:x43:7 vdd x43:nc n046 vdd x43:pfet l=0.6u w=6u
m:x43:8 vdd x43:nb x43:n001 vdd x43:pfet l=0.6u w=6u
m:x43:9 x43:n001 x43:na n046 vdd x43:pfet l=0.6u w=6u
m:x43:10 n046 x43:na x43:n004 0 x43:nfet l=0.6u w=3u
m:x43:11 n046 x43:nb x43:n004 0 x43:nfet l=0.6u w=3u
m:x43:12 x43:n004 x43:nc 0 0 x43:nfet l=0.6u w=3u
m:x43:13 x43:n003 n031 0 0 x43:nfet l=0.6u w=3u
m:x43:14 x43:n002 n020 x43:n003 0 x43:nfet l=0.6u w=3u
m:x43:15 vdd n031 x43:n002 vdd x43:pfet l=0.6u w=3u
m:x43:16 vdd n020 x43:n002 vdd x43:pfet l=0.6u w=3u
m:x43:17 vdd x43:n002 n047 vdd x43:pfet l=0.6u w=3u
m:x43:18 n047 x43:n002 0 0 x43:nfet l=0.6u w=1.5u
m:x44:1 vdd n025 x44:nb vdd x44:pfet l=0.6u w=3u
m:x44:2 x44:nb n025 0 0 x44:nfet l=0.6u w=1.5u
m:x44:3 vdd n034 x44:na vdd x44:pfet l=0.6u w=3u
m:x44:4 x44:na n034 0 0 x44:nfet l=0.6u w=1.5u
m:x44:5 vdd n022 x44:nc vdd x44:pfet l=0.6u w=3u
m:x44:6 x44:nc n022 0 0 x44:nfet l=0.6u w=1.5u
m:x44:7 vdd x44:nc n061 vdd x44:pfet l=0.6u w=6u
m:x44:8 vdd x44:nb x44:n001 vdd x44:pfet l=0.6u w=6u
m:x44:9 x44:n001 x44:na n061 vdd x44:pfet l=0.6u w=6u
m:x44:10 n061 x44:na x44:n004 0 x44:nfet l=0.6u w=3u
m:x44:11 n061 x44:nb x44:n004 0 x44:nfet l=0.6u w=3u
m:x44:12 x44:n004 x44:nc 0 0 x44:nfet l=0.6u w=3u
m:x44:13 x44:n003 n025 0 0 x44:nfet l=0.6u w=3u
m:x44:14 x44:n002 n037 x44:n003 0 x44:nfet l=0.6u w=3u
m:x44:15 vdd n025 x44:n002 vdd x44:pfet l=0.6u w=3u
m:x44:16 vdd n037 x44:n002 vdd x44:pfet l=0.6u w=3u
m:x44:17 vdd x44:n002 n063 vdd x44:pfet l=0.6u w=3u
m:x44:18 n063 x44:n002 0 0 x44:nfet l=0.6u w=1.5u
m:x45:1 vdd n019 x45:nb vdd x45:pfet l=0.6u w=3u
m:x45:2 x45:nb n019 0 0 x45:nfet l=0.6u w=1.5u
m:x45:3 vdd n028 x45:na vdd x45:pfet l=0.6u w=3u
m:x45:4 x45:na n028 0 0 x45:nfet l=0.6u w=1.5u
m:x45:5 vdd n016 x45:nc vdd x45:pfet l=0.6u w=3u
m:x45:6 x45:nc n016 0 0 x45:nfet l=0.6u w=1.5u
m:x45:7 vdd x45:nc n071 vdd x45:pfet l=0.6u w=6u
m:x45:8 vdd x45:nb x45:n001 vdd x45:pfet l=0.6u w=6u
m:x45:9 x45:n001 x45:na n071 vdd x45:pfet l=0.6u w=6u
m:x45:10 n071 x45:na x45:n004 0 x45:nfet l=0.6u w=3u
m:x45:11 n071 x45:nb x45:n004 0 x45:nfet l=0.6u w=3u
m:x45:12 x45:n004 x45:nc 0 0 x45:nfet l=0.6u w=3u
m:x45:13 x45:n003 n019 0 0 x45:nfet l=0.6u w=3u
m:x45:14 x45:n002 n031 x45:n003 0 x45:nfet l=0.6u w=3u
m:x45:15 vdd n019 x45:n002 vdd x45:pfet l=0.6u w=3u
m:x45:16 vdd n031 x45:n002 vdd x45:pfet l=0.6u w=3u
m:x45:17 vdd x45:n002 n072 vdd x45:pfet l=0.6u w=3u
m:x45:18 n072 x45:n002 0 0 x45:nfet l=0.6u w=1.5u
m:x46:1 vdd n045 x46:nb vdd x46:pfet l=0.6u w=3u
m:x46:2 x46:nb n045 0 0 x46:nfet l=0.6u w=1.5u
m:x46:3 vdd n022 x46:na vdd x46:pfet l=0.6u w=3u
m:x46:4 x46:na n022 0 0 x46:nfet l=0.6u w=1.5u
m:x46:5 vdd n044 x46:nc vdd x46:pfet l=0.6u w=3u
m:x46:6 x46:nc n044 0 0 x46:nfet l=0.6u w=1.5u
m:x46:7 vdd x46:nc n069 vdd x46:pfet l=0.6u w=6u
m:x46:8 vdd x46:nb x46:n001 vdd x46:pfet l=0.6u w=6u
m:x46:9 x46:n001 x46:na n069 vdd x46:pfet l=0.6u w=6u
m:x46:10 n069 x46:na x46:n004 0 x46:nfet l=0.6u w=3u
m:x46:11 n069 x46:nb x46:n004 0 x46:nfet l=0.6u w=3u
m:x46:12 x46:n004 x46:nc 0 0 x46:nfet l=0.6u w=3u
m:x46:13 x46:n003 n045 0 0 x46:nfet l=0.6u w=3u
m:x46:14 x46:n002 n025 x46:n003 0 x46:nfet l=0.6u w=3u
m:x46:15 vdd n045 x46:n002 vdd x46:pfet l=0.6u w=3u
m:x46:16 vdd n025 x46:n002 vdd x46:pfet l=0.6u w=3u
m:x46:17 vdd x46:n002 n070 vdd x46:pfet l=0.6u w=3u
m:x46:18 n070 x46:n002 0 0 x46:nfet l=0.6u w=1.5u
m:x47:1 vdd n043 x47:nb vdd x47:pfet l=0.6u w=3u
m:x47:2 x47:nb n043 0 0 x47:nfet l=0.6u w=1.5u
m:x47:3 vdd n016 x47:na vdd x47:pfet l=0.6u w=3u
m:x47:4 x47:na n016 0 0 x47:nfet l=0.6u w=1.5u
m:x47:5 vdd n042 x47:nc vdd x47:pfet l=0.6u w=3u
m:x47:6 x47:nc n042 0 0 x47:nfet l=0.6u w=1.5u
m:x47:7 vdd x47:nc n067 vdd x47:pfet l=0.6u w=6u
m:x47:8 vdd x47:nb x47:n001 vdd x47:pfet l=0.6u w=6u
m:x47:9 x47:n001 x47:na n067 vdd x47:pfet l=0.6u w=6u
m:x47:10 n067 x47:na x47:n004 0 x47:nfet l=0.6u w=3u
m:x47:11 n067 x47:nb x47:n004 0 x47:nfet l=0.6u w=3u
m:x47:12 x47:n004 x47:nc 0 0 x47:nfet l=0.6u w=3u
m:x47:13 x47:n003 n043 0 0 x47:nfet l=0.6u w=3u
m:x47:14 x47:n002 n019 x47:n003 0 x47:nfet l=0.6u w=3u
m:x47:15 vdd n043 x47:n002 vdd x47:pfet l=0.6u w=3u
m:x47:16 vdd n019 x47:n002 vdd x47:pfet l=0.6u w=3u
m:x47:17 vdd x47:n002 n068 vdd x47:pfet l=0.6u w=3u
m:x47:18 n068 x47:n002 0 0 x47:nfet l=0.6u w=1.5u
m:x50:1 vdd x50:n001 n107 vdd x50:pfet l=0.6u w=3u
m:x50:2 n107 x50:n001 0 0 x50:nfet l=0.6u w=1.5u
m:x50:3 vdd n057 x50:n001 vdd x50:pfet l=0.6u w=3u
m:x50:4 x50:n001 n057 0 0 x50:nfet l=0.6u w=1.5u
m:x51:1 vdd x51:n001 n075 vdd x51:pfet l=0.6u w=3u
m:x51:2 n075 x51:n001 0 0 x51:nfet l=0.6u w=1.5u
m:x51:3 vdd n054 x51:n001 vdd x51:pfet l=0.6u w=3u
m:x51:4 x51:n001 n054 0 0 x51:nfet l=0.6u w=1.5u
m:x52:1 vdd n064 x52:nb vdd x52:pfet l=0.6u w=3u
m:x52:2 x52:nb n064 0 0 x52:nfet l=0.6u w=1.5u
m:x52:3 vdd n039 x52:na vdd x52:pfet l=0.6u w=3u
m:x52:4 x52:na n039 0 0 x52:nfet l=0.6u w=1.5u
m:x52:5 vdd n062 x52:nc vdd x52:pfet l=0.6u w=3u
m:x52:6 x52:nc n062 0 0 x52:nfet l=0.6u w=1.5u
m:x52:7 vdd x52:nc n093 vdd x52:pfet l=0.6u w=3u
m:x52:8 vdd x52:na x52:n001 vdd x52:pfet l=0.6u w=3u
m:x52:9 x52:n001 x52:nb n093 vdd x52:pfet l=0.6u w=3u
m:x52:10 n093 x52:na x52:n002 0 x52:nfet l=0.6u w=1.5u
m:x52:11 n093 x52:nb x52:n002 0 x52:nfet l=0.6u w=1.5u
m:x52:12 x52:n002 x52:nc 0 0 x52:nfet l=0.6u w=1.5u
m:x53:1 vdd n059 x53:nb vdd x53:pfet l=0.6u w=3u
m:x53:2 x53:nb n059 0 0 x53:nfet l=0.6u w=1.5u
m:x53:3 vdd n060 x53:na vdd x53:pfet l=0.6u w=3u
m:x53:4 x53:na n060 0 0 x53:nfet l=0.6u w=1.5u
m:x53:5 vdd n058 x53:nc vdd x53:pfet l=0.6u w=3u
m:x53:6 x53:nc n058 0 0 x53:nfet l=0.6u w=1.5u
m:x53:7 vdd x53:nc n074 vdd x53:pfet l=0.6u w=3u
m:x53:8 vdd x53:na x53:n001 vdd x53:pfet l=0.6u w=3u
m:x53:9 x53:n001 x53:nb n074 vdd x53:pfet l=0.6u w=3u
m:x53:10 n074 x53:na x53:n002 0 x53:nfet l=0.6u w=1.5u
m:x53:11 n074 x53:nb x53:n002 0 x53:nfet l=0.6u w=1.5u
m:x53:12 x53:n002 x53:nc 0 0 x53:nfet l=0.6u w=1.5u
m:x54:1 vdd n056 x54:nb vdd x54:pfet l=0.6u w=3u
m:x54:2 x54:nb n056 0 0 x54:nfet l=0.6u w=1.5u
m:x54:3 vdd n057 x54:na vdd x54:pfet l=0.6u w=3u
m:x54:4 x54:na n057 0 0 x54:nfet l=0.6u w=1.5u
m:x54:5 vdd n055 x54:nc vdd x54:pfet l=0.6u w=3u
m:x54:6 x54:nc n055 0 0 x54:nfet l=0.6u w=1.5u
m:x54:7 vdd x54:nc n092 vdd x54:pfet l=0.6u w=3u
m:x54:8 vdd x54:na x54:n001 vdd x54:pfet l=0.6u w=3u
m:x54:9 x54:n001 x54:nb n092 vdd x54:pfet l=0.6u w=3u
m:x54:10 n092 x54:na x54:n002 0 x54:nfet l=0.6u w=1.5u
m:x54:11 n092 x54:nb x54:n002 0 x54:nfet l=0.6u w=1.5u
m:x54:12 x54:n002 x54:nc 0 0 x54:nfet l=0.6u w=1.5u
m:x55:1 vdd n053 x55:nb vdd x55:pfet l=0.6u w=3u
m:x55:2 x55:nb n053 0 0 x55:nfet l=0.6u w=1.5u
m:x55:3 vdd n054 x55:na vdd x55:pfet l=0.6u w=3u
m:x55:4 x55:na n054 0 0 x55:nfet l=0.6u w=1.5u
m:x55:5 vdd n052 x55:nc vdd x55:pfet l=0.6u w=3u
m:x55:6 x55:nc n052 0 0 x55:nfet l=0.6u w=1.5u
m:x55:7 vdd x55:nc n073 vdd x55:pfet l=0.6u w=3u
m:x55:8 vdd x55:na x55:n001 vdd x55:pfet l=0.6u w=3u
m:x55:9 x55:n001 x55:nb n073 vdd x55:pfet l=0.6u w=3u
m:x55:10 n073 x55:na x55:n002 0 x55:nfet l=0.6u w=1.5u
m:x55:11 n073 x55:nb x55:n002 0 x55:nfet l=0.6u w=1.5u
m:x55:12 x55:n002 x55:nc 0 0 x55:nfet l=0.6u w=1.5u
m:x16:1 vdd n051 x16:nb vdd x16:pfet l=0.6u w=3u
m:x16:2 x16:nb n051 0 0 x16:nfet l=0.6u w=1.5u
m:x16:3 vdd n062 x16:na vdd x16:pfet l=0.6u w=3u
m:x16:4 x16:na n062 0 0 x16:nfet l=0.6u w=1.5u
m:x16:5 vdd n050 x16:nc vdd x16:pfet l=0.6u w=3u
m:x16:6 x16:nc n050 0 0 x16:nfet l=0.6u w=1.5u
m:x16:7 vdd x16:nc n090 vdd x16:pfet l=0.6u w=6u
m:x16:8 vdd x16:nb x16:n001 vdd x16:pfet l=0.6u w=6u
m:x16:9 x16:n001 x16:na n090 vdd x16:pfet l=0.6u w=6u
m:x16:10 n090 x16:na x16:n004 0 x16:nfet l=0.6u w=3u
m:x16:11 n090 x16:nb x16:n004 0 x16:nfet l=0.6u w=3u
m:x16:12 x16:n004 x16:nc 0 0 x16:nfet l=0.6u w=3u
m:x16:13 x16:n003 n051 0 0 x16:nfet l=0.6u w=3u
m:x16:14 x16:n002 n064 x16:n003 0 x16:nfet l=0.6u w=3u
m:x16:15 vdd n051 x16:n002 vdd x16:pfet l=0.6u w=3u
m:x16:16 vdd n064 x16:n002 vdd x16:pfet l=0.6u w=3u
m:x16:17 vdd x16:n002 n091 vdd x16:pfet l=0.6u w=3u
m:x16:18 n091 x16:n002 0 0 x16:nfet l=0.6u w=1.5u
m:x33:1 vdd n049 x33:nb vdd x33:pfet l=0.6u w=3u
m:x33:2 x33:nb n049 0 0 x33:nfet l=0.6u w=1.5u
m:x33:3 vdd n058 x33:na vdd x33:pfet l=0.6u w=3u
m:x33:4 x33:na n058 0 0 x33:nfet l=0.6u w=1.5u
m:x33:5 vdd n048 x33:nc vdd x33:pfet l=0.6u w=3u
m:x33:6 x33:nc n048 0 0 x33:nfet l=0.6u w=1.5u
m:x33:7 vdd x33:nc n088 vdd x33:pfet l=0.6u w=6u
m:x33:8 vdd x33:nb x33:n001 vdd x33:pfet l=0.6u w=6u
m:x33:9 x33:n001 x33:na n088 vdd x33:pfet l=0.6u w=6u
m:x33:10 n088 x33:na x33:n004 0 x33:nfet l=0.6u w=3u
m:x33:11 n088 x33:nb x33:n004 0 x33:nfet l=0.6u w=3u
m:x33:12 x33:n004 x33:nc 0 0 x33:nfet l=0.6u w=3u
m:x33:13 x33:n003 n049 0 0 x33:nfet l=0.6u w=3u
m:x33:14 x33:n002 n059 x33:n003 0 x33:nfet l=0.6u w=3u
m:x33:15 vdd n049 x33:n002 vdd x33:pfet l=0.6u w=3u
m:x33:16 vdd n059 x33:n002 vdd x33:pfet l=0.6u w=3u
m:x33:17 vdd x33:n002 n089 vdd x33:pfet l=0.6u w=3u
m:x33:18 n089 x33:n002 0 0 x33:nfet l=0.6u w=1.5u
m:x49:1 vdd n047 x49:nb vdd x49:pfet l=0.6u w=3u
m:x49:2 x49:nb n047 0 0 x49:nfet l=0.6u w=1.5u
m:x49:3 vdd n055 x49:na vdd x49:pfet l=0.6u w=3u
m:x49:4 x49:na n055 0 0 x49:nfet l=0.6u w=1.5u
m:x49:5 vdd n046 x49:nc vdd x49:pfet l=0.6u w=3u
m:x49:6 x49:nc n046 0 0 x49:nfet l=0.6u w=1.5u
m:x49:7 vdd x49:nc n086 vdd x49:pfet l=0.6u w=6u
m:x49:8 vdd x49:nb x49:n001 vdd x49:pfet l=0.6u w=6u
m:x49:9 x49:n001 x49:na n086 vdd x49:pfet l=0.6u w=6u
m:x49:10 n086 x49:na x49:n004 0 x49:nfet l=0.6u w=3u
m:x49:11 n086 x49:nb x49:n004 0 x49:nfet l=0.6u w=3u
m:x49:12 x49:n004 x49:nc 0 0 x49:nfet l=0.6u w=3u
m:x49:13 x49:n003 n047 0 0 x49:nfet l=0.6u w=3u
m:x49:14 x49:n002 n056 x49:n003 0 x49:nfet l=0.6u w=3u
m:x49:15 vdd n047 x49:n002 vdd x49:pfet l=0.6u w=3u
m:x49:16 vdd n056 x49:n002 vdd x49:pfet l=0.6u w=3u
m:x49:17 vdd x49:n002 n087 vdd x49:pfet l=0.6u w=3u
m:x49:18 n087 x49:n002 0 0 x49:nfet l=0.6u w=1.5u
m:x56:1 vdd n063 x56:nb vdd x56:pfet l=0.6u w=3u
m:x56:2 x56:nb n063 0 0 x56:nfet l=0.6u w=1.5u
m:x56:3 vdd n052 x56:na vdd x56:pfet l=0.6u w=3u
m:x56:4 x56:na n052 0 0 x56:nfet l=0.6u w=1.5u
m:x56:5 vdd n061 x56:nc vdd x56:pfet l=0.6u w=3u
m:x56:6 x56:nc n061 0 0 x56:nfet l=0.6u w=1.5u
m:x56:7 vdd x56:nc n084 vdd x56:pfet l=0.6u w=6u
m:x56:8 vdd x56:nb x56:n001 vdd x56:pfet l=0.6u w=6u
m:x56:9 x56:n001 x56:na n084 vdd x56:pfet l=0.6u w=6u
m:x56:10 n084 x56:na x56:n004 0 x56:nfet l=0.6u w=3u
m:x56:11 n084 x56:nb x56:n004 0 x56:nfet l=0.6u w=3u
m:x56:12 x56:n004 x56:nc 0 0 x56:nfet l=0.6u w=3u
m:x56:13 x56:n003 n063 0 0 x56:nfet l=0.6u w=3u
m:x56:14 x56:n002 n053 x56:n003 0 x56:nfet l=0.6u w=3u
m:x56:15 vdd n063 x56:n002 vdd x56:pfet l=0.6u w=3u
m:x56:16 vdd n053 x56:n002 vdd x56:pfet l=0.6u w=3u
m:x56:17 vdd x56:n002 n085 vdd x56:pfet l=0.6u w=3u
m:x56:18 n085 x56:n002 0 0 x56:nfet l=0.6u w=1.5u
m:x57:1 vdd n072 x57:nb vdd x57:pfet l=0.6u w=3u
m:x57:2 x57:nb n072 0 0 x57:nfet l=0.6u w=1.5u
m:x57:3 vdd n050 x57:na vdd x57:pfet l=0.6u w=3u
m:x57:4 x57:na n050 0 0 x57:nfet l=0.6u w=1.5u
m:x57:5 vdd n071 x57:nc vdd x57:pfet l=0.6u w=3u
m:x57:6 x57:nc n071 0 0 x57:nfet l=0.6u w=1.5u
m:x57:7 vdd x57:nc n082 vdd x57:pfet l=0.6u w=6u
m:x57:8 vdd x57:nb x57:n001 vdd x57:pfet l=0.6u w=6u
m:x57:9 x57:n001 x57:na n082 vdd x57:pfet l=0.6u w=6u
m:x57:10 n082 x57:na x57:n004 0 x57:nfet l=0.6u w=3u
m:x57:11 n082 x57:nb x57:n004 0 x57:nfet l=0.6u w=3u
m:x57:12 x57:n004 x57:nc 0 0 x57:nfet l=0.6u w=3u
m:x57:13 x57:n003 n072 0 0 x57:nfet l=0.6u w=3u
m:x57:14 x57:n002 n051 x57:n003 0 x57:nfet l=0.6u w=3u
m:x57:15 vdd n072 x57:n002 vdd x57:pfet l=0.6u w=3u
m:x57:16 vdd n051 x57:n002 vdd x57:pfet l=0.6u w=3u
m:x57:17 vdd x57:n002 n083 vdd x57:pfet l=0.6u w=3u
m:x57:18 n083 x57:n002 0 0 x57:nfet l=0.6u w=1.5u
m:x58:1 vdd n070 x58:nb vdd x58:pfet l=0.6u w=3u
m:x58:2 x58:nb n070 0 0 x58:nfet l=0.6u w=1.5u
m:x58:3 vdd n048 x58:na vdd x58:pfet l=0.6u w=3u
m:x58:4 x58:na n048 0 0 x58:nfet l=0.6u w=1.5u
m:x58:5 vdd n069 x58:nc vdd x58:pfet l=0.6u w=3u
m:x58:6 x58:nc n069 0 0 x58:nfet l=0.6u w=1.5u
m:x58:7 vdd x58:nc n080 vdd x58:pfet l=0.6u w=6u
m:x58:8 vdd x58:nb x58:n001 vdd x58:pfet l=0.6u w=6u
m:x58:9 x58:n001 x58:na n080 vdd x58:pfet l=0.6u w=6u
m:x58:10 n080 x58:na x58:n004 0 x58:nfet l=0.6u w=3u
m:x58:11 n080 x58:nb x58:n004 0 x58:nfet l=0.6u w=3u
m:x58:12 x58:n004 x58:nc 0 0 x58:nfet l=0.6u w=3u
m:x58:13 x58:n003 n070 0 0 x58:nfet l=0.6u w=3u
m:x58:14 x58:n002 n049 x58:n003 0 x58:nfet l=0.6u w=3u
m:x58:15 vdd n070 x58:n002 vdd x58:pfet l=0.6u w=3u
m:x58:16 vdd n049 x58:n002 vdd x58:pfet l=0.6u w=3u
m:x58:17 vdd x58:n002 n081 vdd x58:pfet l=0.6u w=3u
m:x58:18 n081 x58:n002 0 0 x58:nfet l=0.6u w=1.5u
m:x59:1 vdd n068 x59:nb vdd x59:pfet l=0.6u w=3u
m:x59:2 x59:nb n068 0 0 x59:nfet l=0.6u w=1.5u
m:x59:3 vdd n046 x59:na vdd x59:pfet l=0.6u w=3u
m:x59:4 x59:na n046 0 0 x59:nfet l=0.6u w=1.5u
m:x59:5 vdd n067 x59:nc vdd x59:pfet l=0.6u w=3u
m:x59:6 x59:nc n067 0 0 x59:nfet l=0.6u w=1.5u
m:x59:7 vdd x59:nc n078 vdd x59:pfet l=0.6u w=6u
m:x59:8 vdd x59:nb x59:n001 vdd x59:pfet l=0.6u w=6u
m:x59:9 x59:n001 x59:na n078 vdd x59:pfet l=0.6u w=6u
m:x59:10 n078 x59:na x59:n004 0 x59:nfet l=0.6u w=3u
m:x59:11 n078 x59:nb x59:n004 0 x59:nfet l=0.6u w=3u
m:x59:12 x59:n004 x59:nc 0 0 x59:nfet l=0.6u w=3u
m:x59:13 x59:n003 n068 0 0 x59:nfet l=0.6u w=3u
m:x59:14 x59:n002 n047 x59:n003 0 x59:nfet l=0.6u w=3u
m:x59:15 vdd n068 x59:n002 vdd x59:pfet l=0.6u w=3u
m:x59:16 vdd n047 x59:n002 vdd x59:pfet l=0.6u w=3u
m:x59:17 vdd x59:n002 n079 vdd x59:pfet l=0.6u w=3u
m:x59:18 n079 x59:n002 0 0 x59:nfet l=0.6u w=1.5u
m:x61:1 vdd x61:n001 n106 vdd x61:pfet l=0.6u w=3u
m:x61:2 n106 x61:n001 0 0 x61:nfet l=0.6u w=1.5u
m:x61:3 vdd n093 x61:n001 vdd x61:pfet l=0.6u w=3u
m:x61:4 x61:n001 n093 0 0 x61:nfet l=0.6u w=1.5u
m:x62:1 vdd x62:n001 n105 vdd x62:pfet l=0.6u w=3u
m:x62:2 n105 x62:n001 0 0 x62:nfet l=0.6u w=1.5u
m:x62:3 vdd n074 x62:n001 vdd x62:pfet l=0.6u w=3u
m:x62:4 x62:n001 n074 0 0 x62:nfet l=0.6u w=1.5u
m:x63:1 vdd x63:n001 n104 vdd x63:pfet l=0.6u w=3u
m:x63:2 n104 x63:n001 0 0 x63:nfet l=0.6u w=1.5u
m:x63:3 vdd n092 x63:n001 vdd x63:pfet l=0.6u w=3u
m:x63:4 x63:n001 n092 0 0 x63:nfet l=0.6u w=1.5u
m:x64:1 vdd x64:n001 n103 vdd x64:pfet l=0.6u w=3u
m:x64:2 n103 x64:n001 0 0 x64:nfet l=0.6u w=1.5u
m:x64:3 vdd n073 x64:n001 vdd x64:pfet l=0.6u w=3u
m:x64:4 x64:n001 n073 0 0 x64:nfet l=0.6u w=1.5u
m:x65:1 vdd n091 x65:nb vdd x65:pfet l=0.6u w=3u
m:x65:2 x65:nb n091 0 0 x65:nfet l=0.6u w=1.5u
m:x65:3 vdd n060 x65:na vdd x65:pfet l=0.6u w=3u
m:x65:4 x65:na n060 0 0 x65:nfet l=0.6u w=1.5u
m:x65:5 vdd n090 x65:nc vdd x65:pfet l=0.6u w=3u
m:x65:6 x65:nc n090 0 0 x65:nfet l=0.6u w=1.5u
m:x65:7 vdd x65:nc n102 vdd x65:pfet l=0.6u w=3u
m:x65:8 vdd x65:na x65:n001 vdd x65:pfet l=0.6u w=3u
m:x65:9 x65:n001 x65:nb n102 vdd x65:pfet l=0.6u w=3u
m:x65:10 n102 x65:na x65:n002 0 x65:nfet l=0.6u w=1.5u
m:x65:11 n102 x65:nb x65:n002 0 x65:nfet l=0.6u w=1.5u
m:x65:12 x65:n002 x65:nc 0 0 x65:nfet l=0.6u w=1.5u
m:x66:1 vdd n089 x66:nb vdd x66:pfet l=0.6u w=3u
m:x66:2 x66:nb n089 0 0 x66:nfet l=0.6u w=1.5u
m:x66:3 vdd n060 x66:na vdd x66:pfet l=0.6u w=3u
m:x66:4 x66:na n060 0 0 x66:nfet l=0.6u w=1.5u
m:x66:5 vdd n088 x66:nc vdd x66:pfet l=0.6u w=3u
m:x66:6 x66:nc n088 0 0 x66:nfet l=0.6u w=1.5u
m:x66:7 vdd x66:nc n101 vdd x66:pfet l=0.6u w=3u
m:x66:8 vdd x66:na x66:n001 vdd x66:pfet l=0.6u w=3u
m:x66:9 x66:n001 x66:nb n101 vdd x66:pfet l=0.6u w=3u
m:x66:10 n101 x66:na x66:n002 0 x66:nfet l=0.6u w=1.5u
m:x66:11 n101 x66:nb x66:n002 0 x66:nfet l=0.6u w=1.5u
m:x66:12 x66:n002 x66:nc 0 0 x66:nfet l=0.6u w=1.5u
m:x67:1 vdd n087 x67:nb vdd x67:pfet l=0.6u w=3u
m:x67:2 x67:nb n087 0 0 x67:nfet l=0.6u w=1.5u
m:x67:3 vdd n075 x67:na vdd x67:pfet l=0.6u w=3u
m:x67:4 x67:na n075 0 0 x67:nfet l=0.6u w=1.5u
m:x67:5 vdd n086 x67:nc vdd x67:pfet l=0.6u w=3u
m:x67:6 x67:nc n086 0 0 x67:nfet l=0.6u w=1.5u
m:x67:7 vdd x67:nc n100 vdd x67:pfet l=0.6u w=3u
m:x67:8 vdd x67:na x67:n001 vdd x67:pfet l=0.6u w=3u
m:x67:9 x67:n001 x67:nb n100 vdd x67:pfet l=0.6u w=3u
m:x67:10 n100 x67:na x67:n002 0 x67:nfet l=0.6u w=1.5u
m:x67:11 n100 x67:nb x67:n002 0 x67:nfet l=0.6u w=1.5u
m:x67:12 x67:n002 x67:nc 0 0 x67:nfet l=0.6u w=1.5u
m:x68:1 vdd n085 x68:nb vdd x68:pfet l=0.6u w=3u
m:x68:2 x68:nb n085 0 0 x68:nfet l=0.6u w=1.5u
m:x68:3 vdd n075 x68:na vdd x68:pfet l=0.6u w=3u
m:x68:4 x68:na n075 0 0 x68:nfet l=0.6u w=1.5u
m:x68:5 vdd n084 x68:nc vdd x68:pfet l=0.6u w=3u
m:x68:6 x68:nc n084 0 0 x68:nfet l=0.6u w=1.5u
m:x68:7 vdd x68:nc n099 vdd x68:pfet l=0.6u w=3u
m:x68:8 vdd x68:na x68:n001 vdd x68:pfet l=0.6u w=3u
m:x68:9 x68:n001 x68:nb n099 vdd x68:pfet l=0.6u w=3u
m:x68:10 n099 x68:na x68:n002 0 x68:nfet l=0.6u w=1.5u
m:x68:11 n099 x68:nb x68:n002 0 x68:nfet l=0.6u w=1.5u
m:x68:12 x68:n002 x68:nc 0 0 x68:nfet l=0.6u w=1.5u
m:x69:1 vdd n083 x69:nb vdd x69:pfet l=0.6u w=3u
m:x69:2 x69:nb n083 0 0 x69:nfet l=0.6u w=1.5u
m:x69:3 vdd n074 x69:na vdd x69:pfet l=0.6u w=3u
m:x69:4 x69:na n074 0 0 x69:nfet l=0.6u w=1.5u
m:x69:5 vdd n082 x69:nc vdd x69:pfet l=0.6u w=3u
m:x69:6 x69:nc n082 0 0 x69:nfet l=0.6u w=1.5u
m:x69:7 vdd x69:nc n098 vdd x69:pfet l=0.6u w=3u
m:x69:8 vdd x69:na x69:n001 vdd x69:pfet l=0.6u w=3u
m:x69:9 x69:n001 x69:nb n098 vdd x69:pfet l=0.6u w=3u
m:x69:10 n098 x69:na x69:n002 0 x69:nfet l=0.6u w=1.5u
m:x69:11 n098 x69:nb x69:n002 0 x69:nfet l=0.6u w=1.5u
m:x69:12 x69:n002 x69:nc 0 0 x69:nfet l=0.6u w=1.5u
m:x70:1 vdd n081 x70:nb vdd x70:pfet l=0.6u w=3u
m:x70:2 x70:nb n081 0 0 x70:nfet l=0.6u w=1.5u
m:x70:3 vdd n074 x70:na vdd x70:pfet l=0.6u w=3u
m:x70:4 x70:na n074 0 0 x70:nfet l=0.6u w=1.5u
m:x70:5 vdd n080 x70:nc vdd x70:pfet l=0.6u w=3u
m:x70:6 x70:nc n080 0 0 x70:nfet l=0.6u w=1.5u
m:x70:7 vdd x70:nc n097 vdd x70:pfet l=0.6u w=3u
m:x70:8 vdd x70:na x70:n001 vdd x70:pfet l=0.6u w=3u
m:x70:9 x70:n001 x70:nb n097 vdd x70:pfet l=0.6u w=3u
m:x70:10 n097 x70:na x70:n002 0 x70:nfet l=0.6u w=1.5u
m:x70:11 n097 x70:nb x70:n002 0 x70:nfet l=0.6u w=1.5u
m:x70:12 x70:n002 x70:nc 0 0 x70:nfet l=0.6u w=1.5u
m:x71:1 vdd n079 x71:nb vdd x71:pfet l=0.6u w=3u
m:x71:2 x71:nb n079 0 0 x71:nfet l=0.6u w=1.5u
m:x71:3 vdd n073 x71:na vdd x71:pfet l=0.6u w=3u
m:x71:4 x71:na n073 0 0 x71:nfet l=0.6u w=1.5u
m:x71:5 vdd n078 x71:nc vdd x71:pfet l=0.6u w=3u
m:x71:6 x71:nc n078 0 0 x71:nfet l=0.6u w=1.5u
m:x71:7 vdd x71:nc n096 vdd x71:pfet l=0.6u w=3u
m:x71:8 vdd x71:na x71:n001 vdd x71:pfet l=0.6u w=3u
m:x71:9 x71:n001 x71:nb n096 vdd x71:pfet l=0.6u w=3u
m:x71:10 n096 x71:na x71:n002 0 x71:nfet l=0.6u w=1.5u
m:x71:11 n096 x71:nb x71:n002 0 x71:nfet l=0.6u w=1.5u
m:x71:12 x71:n002 x71:nc 0 0 x71:nfet l=0.6u w=1.5u
m:x32:1 vdd x32:na x32:n001 vdd x32:pfet l=0.6u w=6u
m:x32:2 x32:n001 n039 s1 vdd x32:pfet l=0.6u w=6u
m:x32:3 vdd p1 x32:n002 vdd x32:pfet l=0.6u w=6u
m:x32:4 x32:n002 x32:nb s1 vdd x32:pfet l=0.6u w=6u
m:x32:5 s1 p1 x32:n003 0 x32:nfet l=0.6u w=3u
m:x32:6 x32:n003 n039 0 0 x32:nfet l=0.6u w=3u
m:x32:7 s1 x32:na x32:n004 0 x32:nfet l=0.6u w=3u
m:x32:8 x32:n004 x32:nb 0 0 x32:nfet l=0.6u w=3u
m:x32:9 vdd n039 x32:nb vdd x32:pfet l=0.6u w=3u
m:x32:10 x32:nb n039 0 0 x32:nfet l=0.6u w=1.5u
m:x32:11 vdd p1 x32:na vdd x32:pfet l=0.6u w=3u
m:x32:12 x32:na p1 0 0 x32:nfet l=0.6u w=1.5u
m:x48:1 vdd x48:na x48:n001 vdd x48:pfet l=0.6u w=6u
m:x48:2 x48:n001 n060 s2 vdd x48:pfet l=0.6u w=6u
m:x48:3 vdd p2 x48:n002 vdd x48:pfet l=0.6u w=6u
m:x48:4 x48:n002 x48:nb s2 vdd x48:pfet l=0.6u w=6u
m:x48:5 s2 p2 x48:n003 0 x48:nfet l=0.6u w=3u
m:x48:6 x48:n003 n060 0 0 x48:nfet l=0.6u w=3u
m:x48:7 s2 x48:na x48:n004 0 x48:nfet l=0.6u w=3u
m:x48:8 x48:n004 x48:nb 0 0 x48:nfet l=0.6u w=3u
m:x48:9 vdd n060 x48:nb vdd x48:pfet l=0.6u w=3u
m:x48:10 x48:nb n060 0 0 x48:nfet l=0.6u w=1.5u
m:x48:11 vdd p2 x48:na vdd x48:pfet l=0.6u w=3u
m:x48:12 x48:na p2 0 0 x48:nfet l=0.6u w=1.5u
m:x60:1 vdd x60:na x60:n001 vdd x60:pfet l=0.6u w=6u
m:x60:2 x60:n001 n107 s3 vdd x60:pfet l=0.6u w=6u
m:x60:3 vdd p3 x60:n002 vdd x60:pfet l=0.6u w=6u
m:x60:4 x60:n002 x60:nb s3 vdd x60:pfet l=0.6u w=6u
m:x60:5 s3 p3 x60:n003 0 x60:nfet l=0.6u w=3u
m:x60:6 x60:n003 n107 0 0 x60:nfet l=0.6u w=3u
m:x60:7 s3 x60:na x60:n004 0 x60:nfet l=0.6u w=3u
m:x60:8 x60:n004 x60:nb 0 0 x60:nfet l=0.6u w=3u
m:x60:9 vdd n107 x60:nb vdd x60:pfet l=0.6u w=3u
m:x60:10 x60:nb n107 0 0 x60:nfet l=0.6u w=1.5u
m:x60:11 vdd p3 x60:na vdd x60:pfet l=0.6u w=3u
m:x60:12 x60:na p3 0 0 x60:nfet l=0.6u w=1.5u
m:x72:1 vdd x72:na x72:n001 vdd x72:pfet l=0.6u w=6u
m:x72:2 x72:n001 n075 s4 vdd x72:pfet l=0.6u w=6u
m:x72:3 vdd p4 x72:n002 vdd x72:pfet l=0.6u w=6u
m:x72:4 x72:n002 x72:nb s4 vdd x72:pfet l=0.6u w=6u
m:x72:5 s4 p4 x72:n003 0 x72:nfet l=0.6u w=3u
m:x72:6 x72:n003 n075 0 0 x72:nfet l=0.6u w=3u
m:x72:7 s4 x72:na x72:n004 0 x72:nfet l=0.6u w=3u
m:x72:8 x72:n004 x72:nb 0 0 x72:nfet l=0.6u w=3u
m:x72:9 vdd n075 x72:nb vdd x72:pfet l=0.6u w=3u
m:x72:10 x72:nb n075 0 0 x72:nfet l=0.6u w=1.5u
m:x72:11 vdd p4 x72:na vdd x72:pfet l=0.6u w=3u
m:x72:12 x72:na p4 0 0 x72:nfet l=0.6u w=1.5u
m:x73:1 vdd x73:na x73:n001 vdd x73:pfet l=0.6u w=6u
m:x73:2 x73:n001 n106 s5 vdd x73:pfet l=0.6u w=6u
m:x73:3 vdd p5 x73:n002 vdd x73:pfet l=0.6u w=6u
m:x73:4 x73:n002 x73:nb s5 vdd x73:pfet l=0.6u w=6u
m:x73:5 s5 p5 x73:n003 0 x73:nfet l=0.6u w=3u
m:x73:6 x73:n003 n106 0 0 x73:nfet l=0.6u w=3u
m:x73:7 s5 x73:na x73:n004 0 x73:nfet l=0.6u w=3u
m:x73:8 x73:n004 x73:nb 0 0 x73:nfet l=0.6u w=3u
m:x73:9 vdd n106 x73:nb vdd x73:pfet l=0.6u w=3u
m:x73:10 x73:nb n106 0 0 x73:nfet l=0.6u w=1.5u
m:x73:11 vdd p5 x73:na vdd x73:pfet l=0.6u w=3u
m:x73:12 x73:na p5 0 0 x73:nfet l=0.6u w=1.5u
m:x74:1 vdd x74:na x74:n001 vdd x74:pfet l=0.6u w=6u
m:x74:2 x74:n001 n105 s6 vdd x74:pfet l=0.6u w=6u
m:x74:3 vdd p6 x74:n002 vdd x74:pfet l=0.6u w=6u
m:x74:4 x74:n002 x74:nb s6 vdd x74:pfet l=0.6u w=6u
m:x74:5 s6 p6 x74:n003 0 x74:nfet l=0.6u w=3u
m:x74:6 x74:n003 n105 0 0 x74:nfet l=0.6u w=3u
m:x74:7 s6 x74:na x74:n004 0 x74:nfet l=0.6u w=3u
m:x74:8 x74:n004 x74:nb 0 0 x74:nfet l=0.6u w=3u
m:x74:9 vdd n105 x74:nb vdd x74:pfet l=0.6u w=3u
m:x74:10 x74:nb n105 0 0 x74:nfet l=0.6u w=1.5u
m:x74:11 vdd p6 x74:na vdd x74:pfet l=0.6u w=3u
m:x74:12 x74:na p6 0 0 x74:nfet l=0.6u w=1.5u
m:x75:1 vdd x75:na x75:n001 vdd x75:pfet l=0.6u w=6u
m:x75:2 x75:n001 n104 s7 vdd x75:pfet l=0.6u w=6u
m:x75:3 vdd p7 x75:n002 vdd x75:pfet l=0.6u w=6u
m:x75:4 x75:n002 x75:nb s7 vdd x75:pfet l=0.6u w=6u
m:x75:5 s7 p7 x75:n003 0 x75:nfet l=0.6u w=3u
m:x75:6 x75:n003 n104 0 0 x75:nfet l=0.6u w=3u
m:x75:7 s7 x75:na x75:n004 0 x75:nfet l=0.6u w=3u
m:x75:8 x75:n004 x75:nb 0 0 x75:nfet l=0.6u w=3u
m:x75:9 vdd n104 x75:nb vdd x75:pfet l=0.6u w=3u
m:x75:10 x75:nb n104 0 0 x75:nfet l=0.6u w=1.5u
m:x75:11 vdd p7 x75:na vdd x75:pfet l=0.6u w=3u
m:x75:12 x75:na p7 0 0 x75:nfet l=0.6u w=1.5u
m:x76:1 vdd x76:na x76:n001 vdd x76:pfet l=0.6u w=6u
m:x76:2 x76:n001 n103 s8 vdd x76:pfet l=0.6u w=6u
m:x76:3 vdd p8 x76:n002 vdd x76:pfet l=0.6u w=6u
m:x76:4 x76:n002 x76:nb s8 vdd x76:pfet l=0.6u w=6u
m:x76:5 s8 p8 x76:n003 0 x76:nfet l=0.6u w=3u
m:x76:6 x76:n003 n103 0 0 x76:nfet l=0.6u w=3u
m:x76:7 s8 x76:na x76:n004 0 x76:nfet l=0.6u w=3u
m:x76:8 x76:n004 x76:nb 0 0 x76:nfet l=0.6u w=3u
m:x76:9 vdd n103 x76:nb vdd x76:pfet l=0.6u w=3u
m:x76:10 x76:nb n103 0 0 x76:nfet l=0.6u w=1.5u
m:x76:11 vdd p8 x76:na vdd x76:pfet l=0.6u w=3u
m:x76:12 x76:na p8 0 0 x76:nfet l=0.6u w=1.5u
m:x77:1 vdd x77:na x77:n001 vdd x77:pfet l=0.6u w=6u
m:x77:2 x77:n001 n102 s9 vdd x77:pfet l=0.6u w=6u
m:x77:3 vdd p9 x77:n002 vdd x77:pfet l=0.6u w=6u
m:x77:4 x77:n002 x77:nb s9 vdd x77:pfet l=0.6u w=6u
m:x77:5 s9 p9 x77:n003 0 x77:nfet l=0.6u w=3u
m:x77:6 x77:n003 n102 0 0 x77:nfet l=0.6u w=3u
m:x77:7 s9 x77:na x77:n004 0 x77:nfet l=0.6u w=3u
m:x77:8 x77:n004 x77:nb 0 0 x77:nfet l=0.6u w=3u
m:x77:9 vdd n102 x77:nb vdd x77:pfet l=0.6u w=3u
m:x77:10 x77:nb n102 0 0 x77:nfet l=0.6u w=1.5u
m:x77:11 vdd p9 x77:na vdd x77:pfet l=0.6u w=3u
m:x77:12 x77:na p9 0 0 x77:nfet l=0.6u w=1.5u
m:x78:1 vdd x78:na x78:n001 vdd x78:pfet l=0.6u w=6u
m:x78:2 x78:n001 n101 s10 vdd x78:pfet l=0.6u w=6u
m:x78:3 vdd p10 x78:n002 vdd x78:pfet l=0.6u w=6u
m:x78:4 x78:n002 x78:nb s10 vdd x78:pfet l=0.6u w=6u
m:x78:5 s10 p10 x78:n003 0 x78:nfet l=0.6u w=3u
m:x78:6 x78:n003 n101 0 0 x78:nfet l=0.6u w=3u
m:x78:7 s10 x78:na x78:n004 0 x78:nfet l=0.6u w=3u
m:x78:8 x78:n004 x78:nb 0 0 x78:nfet l=0.6u w=3u
m:x78:9 vdd n101 x78:nb vdd x78:pfet l=0.6u w=3u
m:x78:10 x78:nb n101 0 0 x78:nfet l=0.6u w=1.5u
m:x78:11 vdd p10 x78:na vdd x78:pfet l=0.6u w=3u
m:x78:12 x78:na p10 0 0 x78:nfet l=0.6u w=1.5u
m:x79:1 vdd x79:na x79:n001 vdd x79:pfet l=0.6u w=6u
m:x79:2 x79:n001 n100 s11 vdd x79:pfet l=0.6u w=6u
m:x79:3 vdd p11 x79:n002 vdd x79:pfet l=0.6u w=6u
m:x79:4 x79:n002 x79:nb s11 vdd x79:pfet l=0.6u w=6u
m:x79:5 s11 p11 x79:n003 0 x79:nfet l=0.6u w=3u
m:x79:6 x79:n003 n100 0 0 x79:nfet l=0.6u w=3u
m:x79:7 s11 x79:na x79:n004 0 x79:nfet l=0.6u w=3u
m:x79:8 x79:n004 x79:nb 0 0 x79:nfet l=0.6u w=3u
m:x79:9 vdd n100 x79:nb vdd x79:pfet l=0.6u w=3u
m:x79:10 x79:nb n100 0 0 x79:nfet l=0.6u w=1.5u
m:x79:11 vdd p11 x79:na vdd x79:pfet l=0.6u w=3u
m:x79:12 x79:na p11 0 0 x79:nfet l=0.6u w=1.5u
m:x80:1 vdd x80:na x80:n001 vdd x80:pfet l=0.6u w=6u
m:x80:2 x80:n001 n099 s12 vdd x80:pfet l=0.6u w=6u
m:x80:3 vdd p12 x80:n002 vdd x80:pfet l=0.6u w=6u
m:x80:4 x80:n002 x80:nb s12 vdd x80:pfet l=0.6u w=6u
m:x80:5 s12 p12 x80:n003 0 x80:nfet l=0.6u w=3u
m:x80:6 x80:n003 n099 0 0 x80:nfet l=0.6u w=3u
m:x80:7 s12 x80:na x80:n004 0 x80:nfet l=0.6u w=3u
m:x80:8 x80:n004 x80:nb 0 0 x80:nfet l=0.6u w=3u
m:x80:9 vdd n099 x80:nb vdd x80:pfet l=0.6u w=3u
m:x80:10 x80:nb n099 0 0 x80:nfet l=0.6u w=1.5u
m:x80:11 vdd p12 x80:na vdd x80:pfet l=0.6u w=3u
m:x80:12 x80:na p12 0 0 x80:nfet l=0.6u w=1.5u
m:x81:1 vdd x81:na x81:n001 vdd x81:pfet l=0.6u w=6u
m:x81:2 x81:n001 n098 s13 vdd x81:pfet l=0.6u w=6u
m:x81:3 vdd p13 x81:n002 vdd x81:pfet l=0.6u w=6u
m:x81:4 x81:n002 x81:nb s13 vdd x81:pfet l=0.6u w=6u
m:x81:5 s13 p13 x81:n003 0 x81:nfet l=0.6u w=3u
m:x81:6 x81:n003 n098 0 0 x81:nfet l=0.6u w=3u
m:x81:7 s13 x81:na x81:n004 0 x81:nfet l=0.6u w=3u
m:x81:8 x81:n004 x81:nb 0 0 x81:nfet l=0.6u w=3u
m:x81:9 vdd n098 x81:nb vdd x81:pfet l=0.6u w=3u
m:x81:10 x81:nb n098 0 0 x81:nfet l=0.6u w=1.5u
m:x81:11 vdd p13 x81:na vdd x81:pfet l=0.6u w=3u
m:x81:12 x81:na p13 0 0 x81:nfet l=0.6u w=1.5u
m:x82:1 vdd x82:na x82:n001 vdd x82:pfet l=0.6u w=6u
m:x82:2 x82:n001 n097 s14 vdd x82:pfet l=0.6u w=6u
m:x82:3 vdd p14 x82:n002 vdd x82:pfet l=0.6u w=6u
m:x82:4 x82:n002 x82:nb s14 vdd x82:pfet l=0.6u w=6u
m:x82:5 s14 p14 x82:n003 0 x82:nfet l=0.6u w=3u
m:x82:6 x82:n003 n097 0 0 x82:nfet l=0.6u w=3u
m:x82:7 s14 x82:na x82:n004 0 x82:nfet l=0.6u w=3u
m:x82:8 x82:n004 x82:nb 0 0 x82:nfet l=0.6u w=3u
m:x82:9 vdd n097 x82:nb vdd x82:pfet l=0.6u w=3u
m:x82:10 x82:nb n097 0 0 x82:nfet l=0.6u w=1.5u
m:x82:11 vdd p14 x82:na vdd x82:pfet l=0.6u w=3u
m:x82:12 x82:na p14 0 0 x82:nfet l=0.6u w=1.5u
m:x83:1 vdd x83:na x83:n001 vdd x83:pfet l=0.6u w=6u
m:x83:2 x83:n001 n096 s15 vdd x83:pfet l=0.6u w=6u
m:x83:3 vdd p15 x83:n002 vdd x83:pfet l=0.6u w=6u
m:x83:4 x83:n002 x83:nb s15 vdd x83:pfet l=0.6u w=6u
m:x83:5 s15 p15 x83:n003 0 x83:nfet l=0.6u w=3u
m:x83:6 x83:n003 n096 0 0 x83:nfet l=0.6u w=3u
m:x83:7 s15 x83:na x83:n004 0 x83:nfet l=0.6u w=3u
m:x83:8 x83:n004 x83:nb 0 0 x83:nfet l=0.6u w=3u
m:x83:9 vdd n096 x83:nb vdd x83:pfet l=0.6u w=3u
m:x83:10 x83:nb n096 0 0 x83:nfet l=0.6u w=1.5u
m:x83:11 vdd p15 x83:na vdd x83:pfet l=0.6u w=3u
m:x83:12 x83:na p15 0 0 x83:nfet l=0.6u w=1.5u
m:x84:1 vdd p16 x84:nb vdd x84:pfet l=0.6u w=3u
m:x84:2 x84:nb p16 0 0 x84:nfet l=0.6u w=1.5u
m:x84:3 vdd n094 x84:na vdd x84:pfet l=0.6u w=3u
m:x84:4 x84:na n094 0 0 x84:nfet l=0.6u w=1.5u
m:x84:5 vdd n095 x84:nc vdd x84:pfet l=0.6u w=3u
m:x84:6 x84:nc n095 0 0 x84:nfet l=0.6u w=1.5u
m:x84:7 vdd x84:nc cout vdd x84:pfet l=0.6u w=3u
m:x84:8 vdd x84:na x84:n001 vdd x84:pfet l=0.6u w=3u
m:x84:9 x84:n001 x84:nb cout vdd x84:pfet l=0.6u w=3u
m:x84:10 cout x84:na x84:n002 0 x84:nfet l=0.6u w=1.5u
m:x84:11 cout x84:nb x84:n002 0 x84:nfet l=0.6u w=1.5u
m:x84:12 x84:n002 x84:nc 0 0 x84:nfet l=0.6u w=1.5u
m:x85:1 vdd p15 x85:nb vdd x85:pfet l=0.6u w=3u
m:x85:2 x85:nb p15 0 0 x85:nfet l=0.6u w=1.5u
m:x85:3 vdd n001 x85:na vdd x85:pfet l=0.6u w=3u
m:x85:4 x85:na n001 0 0 x85:nfet l=0.6u w=1.5u
m:x85:5 vdd n015 x85:nc vdd x85:pfet l=0.6u w=3u
m:x85:6 x85:nc n015 0 0 x85:nfet l=0.6u w=1.5u
m:x85:7 vdd x85:nc n040 vdd x85:pfet l=0.6u w=6u
m:x85:8 vdd x85:nb x85:n001 vdd x85:pfet l=0.6u w=6u
m:x85:9 x85:n001 x85:na n040 vdd x85:pfet l=0.6u w=6u
m:x85:10 n040 x85:na x85:n004 0 x85:nfet l=0.6u w=3u
m:x85:11 n040 x85:nb x85:n004 0 x85:nfet l=0.6u w=3u
m:x85:12 x85:n004 x85:nc 0 0 x85:nfet l=0.6u w=3u
m:x85:13 x85:n003 p15 0 0 x85:nfet l=0.6u w=3u
m:x85:14 x85:n002 p14 x85:n003 0 x85:nfet l=0.6u w=3u
m:x85:15 vdd p15 x85:n002 vdd x85:pfet l=0.6u w=3u
m:x85:16 vdd p14 x85:n002 vdd x85:pfet l=0.6u w=3u
m:x85:17 vdd x85:n002 n041 vdd x85:pfet l=0.6u w=3u
m:x85:18 n041 x85:n002 0 0 x85:nfet l=0.6u w=1.5u
m:x86:1 vdd n041 x86:nb vdd x86:pfet l=0.6u w=3u
m:x86:2 x86:nb n041 0 0 x86:nfet l=0.6u w=1.5u
m:x86:3 vdd n022 x86:na vdd x86:pfet l=0.6u w=3u
m:x86:4 x86:na n022 0 0 x86:nfet l=0.6u w=1.5u
m:x86:5 vdd n040 x86:nc vdd x86:pfet l=0.6u w=3u
m:x86:6 x86:nc n040 0 0 x86:nfet l=0.6u w=1.5u
m:x86:7 vdd x86:nc n065 vdd x86:pfet l=0.6u w=6u
m:x86:8 vdd x86:nb x86:n001 vdd x86:pfet l=0.6u w=6u
m:x86:9 x86:n001 x86:na n065 vdd x86:pfet l=0.6u w=6u
m:x86:10 n065 x86:na x86:n004 0 x86:nfet l=0.6u w=3u
m:x86:11 n065 x86:nb x86:n004 0 x86:nfet l=0.6u w=3u
m:x86:12 x86:n004 x86:nc 0 0 x86:nfet l=0.6u w=3u
m:x86:13 x86:n003 n041 0 0 x86:nfet l=0.6u w=3u
m:x86:14 x86:n002 n025 x86:n003 0 x86:nfet l=0.6u w=3u
m:x86:15 vdd n041 x86:n002 vdd x86:pfet l=0.6u w=3u
m:x86:16 vdd n025 x86:n002 vdd x86:pfet l=0.6u w=3u
m:x86:17 vdd x86:n002 n066 vdd x86:pfet l=0.6u w=3u
m:x86:18 n066 x86:n002 0 0 x86:nfet l=0.6u w=1.5u
m:x87:1 vdd n066 x87:nb vdd x87:pfet l=0.6u w=3u
m:x87:2 x87:nb n066 0 0 x87:nfet l=0.6u w=1.5u
m:x87:3 vdd n061 x87:na vdd x87:pfet l=0.6u w=3u
m:x87:4 x87:na n061 0 0 x87:nfet l=0.6u w=1.5u
m:x87:5 vdd n065 x87:nc vdd x87:pfet l=0.6u w=3u
m:x87:6 x87:nc n065 0 0 x87:nfet l=0.6u w=1.5u
m:x87:7 vdd x87:nc n076 vdd x87:pfet l=0.6u w=6u
m:x87:8 vdd x87:nb x87:n001 vdd x87:pfet l=0.6u w=6u
m:x87:9 x87:n001 x87:na n076 vdd x87:pfet l=0.6u w=6u
m:x87:10 n076 x87:na x87:n004 0 x87:nfet l=0.6u w=3u
m:x87:11 n076 x87:nb x87:n004 0 x87:nfet l=0.6u w=3u
m:x87:12 x87:n004 x87:nc 0 0 x87:nfet l=0.6u w=3u
m:x87:13 x87:n003 n066 0 0 x87:nfet l=0.6u w=3u
m:x87:14 x87:n002 n063 x87:n003 0 x87:nfet l=0.6u w=3u
m:x87:15 vdd n066 x87:n002 vdd x87:pfet l=0.6u w=3u
m:x87:16 vdd n063 x87:n002 vdd x87:pfet l=0.6u w=3u
m:x87:17 vdd x87:n002 n077 vdd x87:pfet l=0.6u w=3u
m:x87:18 n077 x87:n002 0 0 x87:nfet l=0.6u w=1.5u
m:x88:1 vdd n077 x88:nb vdd x88:pfet l=0.6u w=3u
m:x88:2 x88:nb n077 0 0 x88:nfet l=0.6u w=1.5u
m:x88:3 vdd n073 x88:na vdd x88:pfet l=0.6u w=3u
m:x88:4 x88:na n073 0 0 x88:nfet l=0.6u w=1.5u
m:x88:5 vdd n076 x88:nc vdd x88:pfet l=0.6u w=3u
m:x88:6 x88:nc n076 0 0 x88:nfet l=0.6u w=1.5u
m:x88:7 vdd x88:nc n094 vdd x88:pfet l=0.6u w=3u
m:x88:8 vdd x88:na x88:n001 vdd x88:pfet l=0.6u w=3u
m:x88:9 x88:n001 x88:nb n094 vdd x88:pfet l=0.6u w=3u
m:x88:10 n094 x88:na x88:n002 0 x88:nfet l=0.6u w=1.5u
m:x88:11 n094 x88:nb x88:n002 0 x88:nfet l=0.6u w=1.5u
m:x88:12 x88:n002 x88:nc 0 0 x88:nfet l=0.6u w=1.5u
m:x89:1 vdd x89:na x89:n001 vdd x89:pfet l=0.6u w=6u
m:x89:2 x89:n001 b16 p16 vdd x89:pfet l=0.6u w=6u
m:x89:3 vdd a16 x89:n002 vdd x89:pfet l=0.6u w=6u
m:x89:4 x89:n002 x89:nb p16 vdd x89:pfet l=0.6u w=6u
m:x89:5 p16 b16 x89:n004 0 x89:nfet l=0.6u w=3u
m:x89:6 x89:n004 a16 0 0 x89:nfet l=0.6u w=3u
m:x89:7 p16 x89:nb x89:n005 0 x89:nfet l=0.6u w=3u
m:x89:8 x89:n005 x89:na 0 0 x89:nfet l=0.6u w=3u
m:x89:9 vdd b16 x89:nb vdd x89:pfet l=0.6u w=3u
m:x89:10 x89:nb b16 0 0 x89:nfet l=0.6u w=1.5u
m:x89:11 vdd a16 x89:na vdd x89:pfet l=0.6u w=3u
m:x89:12 x89:na a16 0 0 x89:nfet l=0.6u w=1.5u
m:x89:13 x89:nand b16 x89:n003 0 x89:nfet l=0.6u w=3u
m:x89:14 x89:n003 a16 0 0 x89:nfet l=0.6u w=3u
m:x89:15 vdd a16 x89:nand vdd x89:pfet l=0.6u w=3u
m:x89:16 vdd b16 x89:nand vdd x89:pfet l=0.6u w=3u
m:x89:17 vdd x89:nand n095 vdd x89:pfet l=0.6u w=3u
m:x89:18 n095 x89:nand 0 0 x89:nfet l=0.6u w=1.5u
m:x90:1 vdd x90:na x90:n001 vdd x90:pfet l=0.6u w=6u
m:x90:2 x90:n001 n094 s16 vdd x90:pfet l=0.6u w=6u
m:x90:3 vdd p16 x90:n002 vdd x90:pfet l=0.6u w=6u
m:x90:4 x90:n002 x90:nb s16 vdd x90:pfet l=0.6u w=6u
m:x90:5 s16 p16 x90:n003 0 x90:nfet l=0.6u w=3u
m:x90:6 x90:n003 n094 0 0 x90:nfet l=0.6u w=3u
m:x90:7 s16 x90:na x90:n004 0 x90:nfet l=0.6u w=3u
m:x90:8 x90:n004 x90:nb 0 0 x90:nfet l=0.6u w=3u
m:x90:9 vdd n094 x90:nb vdd x90:pfet l=0.6u w=3u
m:x90:10 x90:nb n094 0 0 x90:nfet l=0.6u w=1.5u
m:x90:11 vdd p16 x90:na vdd x90:pfet l=0.6u w=3u
.model x90:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x90:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x89:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x89:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x88:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x88:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x87:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x87:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x86:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x86:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x85:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x85:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x84:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x84:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x83:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x83:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x82:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x82:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x81:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x81:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x80:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x80:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x79:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x79:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x78:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x78:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x77:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x77:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x76:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x76:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x75:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x75:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x74:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x74:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x73:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x73:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x72:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x72:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x60:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x60:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x48:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x48:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x32:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x32:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x71:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x71:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x70:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x70:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x69:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x69:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x68:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x68:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x67:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x67:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x66:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x66:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x65:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x65:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x64:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x64:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x63:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x63:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x62:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x62:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x61:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x61:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x59:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x59:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x58:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x58:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x57:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x57:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x56:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x56:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x49:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x49:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x33:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x33:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x16:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x16:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x55:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x55:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x54:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x54:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x53:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x53:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x52:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x52:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x51:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x51:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x50:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x50:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x47:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x47:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x46:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x46:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x45:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x45:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x44:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x44:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x43:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x43:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x42:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x42:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x41:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x41:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x40:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x40:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x39:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x39:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x38:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x38:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x37:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x37:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x36:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x36:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x35:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x35:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x34:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x34:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x31:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x31:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x30:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x30:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x29:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x29:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x28:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x28:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x27:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x27:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x26:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x26:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x25:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x25:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x24:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x24:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x23:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x23:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x22:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x22:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x21:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x21:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x20:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x20:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x19:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x19:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x18:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x18:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x17:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x17:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x15:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x15:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x14:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x14:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x13:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x13:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x12:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x12:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x11:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x11:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x10:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x10:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x9:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x9:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x8:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x8:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x7:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x7:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x6:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x6:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x5:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x5:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x4:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x4:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x3:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x3:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x2:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x2:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
.model x1:pfet pmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=-0.9179952 k1=0.5575604 k2=0.010265 k3=14.0655075 k3b=-2.3032921 w0=1.147829e-6 nlx=1.114768e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=2.2896412 dvt1=0.5213085 dvt2=-0.1337987 u0=202.4540953 ua=2.290194e-9 ub=9.779742e-19 uc=-3.69771e-11 vsat=1.307891e5 a0=0.8356881 ags=0.1568774 b0=2.365956e-6 b1=5e-6 keta=-5.769328e-3 a1=0 a2=1 rdsw=2.746814e3 prwg=2.34865e-3 prwb=0.0172298 wr=1 wint=2.586255e-7 lint=7.205014e-8 xl=0 xw=0 dwg=-2.133054e-8 dwb=9.857534e-9 voff=-0.0837499 nfactor=1.2415529 cit=0 cdsc=4.363744e-4 cdscd=0 cdscb=0 eta0=0.11276 etab=-2.9484e-3 dsub=0.3389402 pclm=4.9847806 pdiblc1=2.481735e-5 pdiblc2=0.01 pdiblcb=0 drout=0.9975107 pscbe1=3.497872e9 pscbe2=4.974352e-9 pvag=10.9914549 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=2.4e-10 cgso=2.4e-10 cgbo=0 cj=7.273568e-4 pb=0.9665597 mj=0.4959837 cjsw=3.114708e-10 pbsw=0.99 mjsw=0.2653654 pvth0=9.420541e-3 prdsw=-231.2571566 pk2=1.396684e-3 wketa=1.862966e-3 lketa=5.728589e-3)
.model x1:nfet nmos (level=49 version=3.1 tnom=27 tox=1.41e-8 xj=1.5e-7 nch=1.7e17 vth0=0.7086 k1=0.8354582 k2=-0.088431 k3=41.4403818 k3b=-14 w0=6.480766e-7 nlx=1e-10 dvt0w=0 dvt1w=5.3e6 dvt2w=-0.032 dvt0=3.6139113 dvt1=0.3795745 dvt2=-0.1399976 u0=533.6953445 ua=7.558023e-10 ub=1.181167e-18 uc=2.582756e-11 vsat=1.300981e5 a0=0.5292985 ags=0.1463715 b0=1.283336e-6 b1=1.408099e-6 keta=-0.0173166 a1=0 a2=1 rdsw=2.268366e3 prwg=-1e-3 prwb=6.320549e-5 wr=1 wint=2.043512e-7 lint=3.034496e-8 xl=0 xw=0 dwg=-1.446149e-8 dwb=2.077539e-8 voff=-0.1137226 nfactor=1.2880596 cit=0 cdsc=1.506004e-4 cdscd=0 cdscb=0 eta0=3.815372e-4 etab=-1.029178e-3 dsub=2.173055e-4 pclm=0.6171774 pdiblc1=0.185986 pdiblc2=3.473187e-3 pdiblcb=-1e-3 drout=0.4037723 pscbe1=5.998012e9 pscbe2=3.788068e-8 pvag=0.012927 delta=0.01 mobmod=1 prt=0 ute=-1.5 kt1=-0.11 kt1l=0 kt2=0.022 ua1=4.31e-9 ub1=-7.61e-18 uc1=-5.6e-11 at=3.3e4 wl=0 wln=1 ww=0 wwn=1 wwl=0 ll=0 lln=1 lw=0 lwn=1 lwl=0 capmod=2 xpart=0.4 cgdo=1.99e-10 cgso=1.99e-10 cgbo=0 cj=4.233802e-4 pb=0.9899238 mj=0.4495859 cjsw=3.825632e-10 pbsw=0.1082556 mjsw=0.1083618 pvth0=0.0212852 prdsw=-16.1546703 pk2=0.0253069 wketa=0.0188633 lketa=0.0204965)
m:x90:12 x90:na p16 0 0 x90:nfet l=0.6u w=1.5u
.end
